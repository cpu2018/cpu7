`default_nettype none

module floor(
  input wire [31:0] x1,
  output wire [31:0] y );

  wire s1, s;
  wire [7:0] e1, e;
  wire [22:0] m1, m;
  assign s1 = x1[31:31];
  assign e1 = x1[30:23];
  assign m1 = x1[22:0];

  wire [24:0] m_25;
  assign m_25 = (e1 >= 8'b10010110) ? {2'b01, m1} :

                ({s1, e1} == 9'b010010101) ? {2'b01, m1[22:1], 1'b0} :
                ({s1, e1} == 9'b010010100) ? {2'b01, m1[22:2], 2'b0} :
                ({s1, e1} == 9'b010010011) ? {2'b01, m1[22:3], 3'b0} :
                ({s1, e1} == 9'b010010010) ? {2'b01, m1[22:4], 4'b0} :
                ({s1, e1} == 9'b010010001) ? {2'b01, m1[22:5], 5'b0} :
                ({s1, e1} == 9'b010010000) ? {2'b01, m1[22:6], 6'b0} :
                ({s1, e1} == 9'b010001111) ? {2'b01, m1[22:7], 7'b0} :
                ({s1, e1} == 9'b010001110) ? {2'b01, m1[22:8], 8'b0} :
                ({s1, e1} == 9'b010001101) ? {2'b01, m1[22:9], 9'b0} :
                ({s1, e1} == 9'b010001100) ? {2'b01, m1[22:10], 10'b0} :
                ({s1, e1} == 9'b010001011) ? {2'b01, m1[22:11], 11'b0} :
                ({s1, e1} == 9'b010001010) ? {2'b01, m1[22:12], 12'b0} :
                ({s1, e1} == 9'b010001001) ? {2'b01, m1[22:13], 13'b0} :
                ({s1, e1} == 9'b010001000) ? {2'b01, m1[22:14], 14'b0} :
                ({s1, e1} == 9'b010000111) ? {2'b01, m1[22:15], 15'b0} :
                ({s1, e1} == 9'b010000110) ? {2'b01, m1[22:16], 16'b0} :
                ({s1, e1} == 9'b010000101) ? {2'b01, m1[22:17], 17'b0} :
                ({s1, e1} == 9'b010000100) ? {2'b01, m1[22:18], 18'b0} :
                ({s1, e1} == 9'b010000011) ? {2'b01, m1[22:19], 19'b0} :
                ({s1, e1} == 9'b010000010) ? {2'b01, m1[22:20], 20'b0} :
                ({s1, e1} == 9'b010000001) ? {2'b01, m1[22:21], 21'b0} :
                ({s1, e1} == 9'b010000000) ? {2'b01, m1[22:22], 22'b0} :
                ({s1, e1} == 9'b001111111) ? {2'b01, 23'b0} :

                ({s1, e1} == 9'b110010101) ? {2'b01, m1[22:1], 1'b0} + {23'b0, m1[0:0], 1'b0} :
                ({s1, e1} == 9'b110010100) ? {2'b01, m1[22:2], 2'b0} + {22'b0, |(m1[1:0]), 2'b0} :
                ({s1, e1} == 9'b110010011) ? {2'b01, m1[22:3], 3'b0} + {21'b0, |(m1[2:0]), 3'b0} :
                ({s1, e1} == 9'b110010010) ? {2'b01, m1[22:4], 4'b0} + {20'b0, |(m1[3:0]), 4'b0} :
                ({s1, e1} == 9'b110010001) ? {2'b01, m1[22:5], 5'b0} + {19'b0, |(m1[4:0]), 5'b0} :
                ({s1, e1} == 9'b110010000) ? {2'b01, m1[22:6], 6'b0} + {18'b0, |(m1[5:0]), 6'b0} :
                ({s1, e1} == 9'b110001111) ? {2'b01, m1[22:7], 7'b0} + {17'b0, |(m1[6:0]), 7'b0} :
                ({s1, e1} == 9'b110001110) ? {2'b01, m1[22:8], 8'b0} + {16'b0, |(m1[7:0]), 8'b0} :
                ({s1, e1} == 9'b110001101) ? {2'b01, m1[22:9], 9'b0} + {15'b0, |(m1[8:0]), 9'b0} :
                ({s1, e1} == 9'b110001100) ? {2'b01, m1[22:10], 10'b0} + {14'b0, |(m1[9:0]), 10'b0} :
                ({s1, e1} == 9'b110001011) ? {2'b01, m1[22:11], 11'b0} + {13'b0, |(m1[10:0]), 11'b0} :
                ({s1, e1} == 9'b110001010) ? {2'b01, m1[22:12], 12'b0} + {12'b0, |(m1[11:0]), 12'b0} :
                ({s1, e1} == 9'b110001001) ? {2'b01, m1[22:13], 13'b0} + {11'b0, |(m1[12:0]), 13'b0} :
                ({s1, e1} == 9'b110001000) ? {2'b01, m1[22:14], 14'b0} + {10'b0, |(m1[13:0]), 14'b0} :
                ({s1, e1} == 9'b110000111) ? {2'b01, m1[22:15], 15'b0} + {9'b0, |(m1[14:0]), 15'b0} :
                ({s1, e1} == 9'b110000110) ? {2'b01, m1[22:16], 16'b0} + {8'b0, |(m1[15:0]), 16'b0} :
                ({s1, e1} == 9'b110000101) ? {2'b01, m1[22:17], 17'b0} + {7'b0, |(m1[16:0]), 17'b0} :
                ({s1, e1} == 9'b110000100) ? {2'b01, m1[22:18], 18'b0} + {6'b0, |(m1[17:0]), 18'b0} :
                ({s1, e1} == 9'b110000011) ? {2'b01, m1[22:19], 19'b0} + {5'b0, |(m1[18:0]), 19'b0} :
                ({s1, e1} == 9'b110000010) ? {2'b01, m1[22:20], 20'b0} + {4'b0, |(m1[19:0]), 20'b0} :
                ({s1, e1} == 9'b110000001) ? {2'b01, m1[22:21], 21'b0} + {3'b0, |(m1[20:0]), 21'b0} :
                ({s1, e1} == 9'b110000000) ? {2'b01, m1[22:22], 22'b0} + {2'b0, |(m1[21:0]), 22'b0} :
                ({s1, e1} == 9'b101111111) ? {2'b01, 23'b0} + {1'b0, |(m1[22:0]), 23'b0} :

                (s1 && {e1, m1} != 31'b0) ? {1'b1, 23'b0, 1'b1} : 25'b0;

  assign s = s1;
  assign e = (m_25[24:24] && m_25[0:0]) ? 8'b01111111 :
             (m_25[24:24]) ? e1 + 8'b1 :
             (m_25[23:23]) ? e1 : 8'b0;
  assign m = (m_25[24:24]) ? m_25[23:1] : m_25[22:0];
  assign y = {s, e, m};

endmodule

`default_nettype wire
