`default_nettype none

module ftoi(
  input wire [31:0] f,
  output wire [31:0] i );

  wire s;
  wire [7:0] e;
  wire [22:0] m;
  assign s = f[31:31];
  assign e = f[30:23];
  assign m = f[22:0];

  wire [23:0] ui24;
  wire [31:0] ui32;
  wire [32:0] uineg33;
  assign ui24 = {1'b1, m};
  assign ui32 = (f == 32'b11001111000000000000000000000000) ? {1'b1, 31'b0} :
                (e >= 8'b10011110) ? 32'b01111111111111111111111111111111 :
                (e == 8'b10011101) ? {1'b0, ui24, 7'b0} :
                (e == 8'b10011100) ? {2'b0, ui24, 6'b0} :
                (e == 8'b10011011) ? {3'b0, ui24, 5'b0} :
                (e == 8'b10011010) ? {4'b0, ui24, 4'b0} :
                (e == 8'b10011001) ? {5'b0, ui24, 3'b0} :
                (e == 8'b10011000) ? {6'b0, ui24, 2'b0} :
                (e == 8'b10010111) ? {7'b0, ui24, 1'b0} :
                (e == 8'b10010110) ? {8'b0, ui24} :
                (e == 8'b10010101) ? {9'b0, ui24[23:1]} + {31'b0, ui24[0:0]} :
                (e == 8'b10010100) ? {10'b0, ui24[23:2]} + {31'b0, ui24[1:1]} :
                (e == 8'b10010011) ? {11'b0, ui24[23:3]} + {31'b0, ui24[2:2]} :
                (e == 8'b10010010) ? {12'b0, ui24[23:4]} + {31'b0, ui24[3:3]} :
                (e == 8'b10010001) ? {13'b0, ui24[23:5]} + {31'b0, ui24[4:4]} :
                (e == 8'b10010000) ? {14'b0, ui24[23:6]} + {31'b0, ui24[5:5]} :
                (e == 8'b10001111) ? {15'b0, ui24[23:7]} + {31'b0, ui24[6:6]} :
                (e == 8'b10001110) ? {16'b0, ui24[23:8]} + {31'b0, ui24[7:7]} :
                (e == 8'b10001101) ? {17'b0, ui24[23:9]} + {31'b0, ui24[8:8]} :
                (e == 8'b10001100) ? {18'b0, ui24[23:10]} + {31'b0, ui24[9:9]} :
                (e == 8'b10001011) ? {19'b0, ui24[23:11]} + {31'b0, ui24[10:10]} :
                (e == 8'b10001010) ? {20'b0, ui24[23:12]} + {31'b0, ui24[11:11]} :
                (e == 8'b10001001) ? {21'b0, ui24[23:13]} + {31'b0, ui24[12:12]} :
                (e == 8'b10001000) ? {22'b0, ui24[23:14]} + {31'b0, ui24[13:13]} :
                (e == 8'b10000111) ? {23'b0, ui24[23:15]} + {31'b0, ui24[14:14]} :
                (e == 8'b10000110) ? {24'b0, ui24[23:16]} + {31'b0, ui24[15:15]} :
                (e == 8'b10000101) ? {25'b0, ui24[23:17]} + {31'b0, ui24[16:16]} :
                (e == 8'b10000100) ? {26'b0, ui24[23:18]} + {31'b0, ui24[17:17]} :
                (e == 8'b10000011) ? {27'b0, ui24[23:19]} + {31'b0, ui24[18:18]} :
                (e == 8'b10000010) ? {28'b0, ui24[23:20]} + {31'b0, ui24[19:19]} :
                (e == 8'b10000001) ? {29'b0, ui24[23:21]} + {31'b0, ui24[20:20]} :
                (e == 8'b10000000) ? {30'b0, ui24[23:22]} + {31'b0, ui24[21:21]} :
                (e == 8'b01111111) ? {31'b0, ui24[23:23]} + {31'b0, ui24[22:22]} :
                (e == 8'b01111110) ? 32'b1 : 32'b0;

assign uineg33 = {1'b0, ~ui32} + 33'b1;

assign i = (ui32 == 32'b0 || ~s) ? ui32 : uineg33[31:0];

endmodule

`default_nettype wire
