`default_nettype none

module fsqrt0(
  input wire [31:0] x1,
  output wire [23:0] y1,
  output wire [23:0] y2 );
  
  function [22:0] fsqrt_table (
    input [9:0] e_m );
    begin
      case(e_m)

10'b0000000000: fsqrt_table = 23'b01101010000010011110011;
10'b0000000001: fsqrt_table = 23'b01101010011001000101111;
10'b0000000010: fsqrt_table = 23'b01101010101111101011111;
10'b0000000011: fsqrt_table = 23'b01101011000110010000100;
10'b0000000100: fsqrt_table = 23'b01101011011100110011110;
10'b0000000101: fsqrt_table = 23'b01101011110011010101101;
10'b0000000110: fsqrt_table = 23'b01101100001001110110000;
10'b0000000111: fsqrt_table = 23'b01101100100000010101001;
10'b0000001000: fsqrt_table = 23'b01101100110110110010110;
10'b0000001001: fsqrt_table = 23'b01101101001101001111000;
10'b0000001010: fsqrt_table = 23'b01101101100011101001111;
10'b0000001011: fsqrt_table = 23'b01101101111010000011100;
10'b0000001100: fsqrt_table = 23'b01101110010000011011101;
10'b0000001101: fsqrt_table = 23'b01101110100110110010011;
10'b0000001110: fsqrt_table = 23'b01101110111101000111111;
10'b0000001111: fsqrt_table = 23'b01101111010011011011111;
10'b0000010000: fsqrt_table = 23'b01101111101001101110101;
10'b0000010001: fsqrt_table = 23'b01110000000000000000000;
10'b0000010010: fsqrt_table = 23'b01110000010110010000000;
10'b0000010011: fsqrt_table = 23'b01110000101100011110110;
10'b0000010100: fsqrt_table = 23'b01110001000010101100000;
10'b0000010101: fsqrt_table = 23'b01110001011000111000000;
10'b0000010110: fsqrt_table = 23'b01110001101111000010110;
10'b0000010111: fsqrt_table = 23'b01110010000101001100001;
10'b0000011000: fsqrt_table = 23'b01110010011011010100001;
10'b0000011001: fsqrt_table = 23'b01110010110001011010110;
10'b0000011010: fsqrt_table = 23'b01110011000111100000001;
10'b0000011011: fsqrt_table = 23'b01110011011101100100010;
10'b0000011100: fsqrt_table = 23'b01110011110011100111000;
10'b0000011101: fsqrt_table = 23'b01110100001001101000100;
10'b0000011110: fsqrt_table = 23'b01110100011111101000101;
10'b0000011111: fsqrt_table = 23'b01110100110101100111100;
10'b0000100000: fsqrt_table = 23'b01110101001011100101000;
10'b0000100001: fsqrt_table = 23'b01110101100001100001011;
10'b0000100010: fsqrt_table = 23'b01110101110111011100010;
10'b0000100011: fsqrt_table = 23'b01110110001101010110000;
10'b0000100100: fsqrt_table = 23'b01110110100011001110011;
10'b0000100101: fsqrt_table = 23'b01110110111001000101101;
10'b0000100110: fsqrt_table = 23'b01110111001110111011011;
10'b0000100111: fsqrt_table = 23'b01110111100100110000000;
10'b0000101000: fsqrt_table = 23'b01110111111010100011011;
10'b0000101001: fsqrt_table = 23'b01111000010000010101011;
10'b0000101010: fsqrt_table = 23'b01111000100110000110010;
10'b0000101011: fsqrt_table = 23'b01111000111011110101110;
10'b0000101100: fsqrt_table = 23'b01111001010001100100001;
10'b0000101101: fsqrt_table = 23'b01111001100111010001001;
10'b0000101110: fsqrt_table = 23'b01111001111100111101000;
10'b0000101111: fsqrt_table = 23'b01111010010010100111100;
10'b0000110000: fsqrt_table = 23'b01111010101000010000111;
10'b0000110001: fsqrt_table = 23'b01111010111101111000111;
10'b0000110010: fsqrt_table = 23'b01111011010011011111110;
10'b0000110011: fsqrt_table = 23'b01111011101001000101011;
10'b0000110100: fsqrt_table = 23'b01111011111110101001110;
10'b0000110101: fsqrt_table = 23'b01111100010100001100111;
10'b0000110110: fsqrt_table = 23'b01111100101001101110111;
10'b0000110111: fsqrt_table = 23'b01111100111111001111101;
10'b0000111000: fsqrt_table = 23'b01111101010100101111001;
10'b0000111001: fsqrt_table = 23'b01111101101010001101100;
10'b0000111010: fsqrt_table = 23'b01111101111111101010100;
10'b0000111011: fsqrt_table = 23'b01111110010101000110100;
10'b0000111100: fsqrt_table = 23'b01111110101010100001001;
10'b0000111101: fsqrt_table = 23'b01111110111111111010101;
10'b0000111110: fsqrt_table = 23'b01111111010101010011000;
10'b0000111111: fsqrt_table = 23'b01111111101010101010001;
10'b0001000000: fsqrt_table = 23'b10000000000000000000000;
10'b0001000001: fsqrt_table = 23'b10000000010101010100110;
10'b0001000010: fsqrt_table = 23'b10000000101010101000010;
10'b0001000011: fsqrt_table = 23'b10000000111111111010101;
10'b0001000100: fsqrt_table = 23'b10000001010101001011111;
10'b0001000101: fsqrt_table = 23'b10000001101010011011111;
10'b0001000110: fsqrt_table = 23'b10000001111111101010110;
10'b0001000111: fsqrt_table = 23'b10000010010100111000100;
10'b0001001000: fsqrt_table = 23'b10000010101010000101000;
10'b0001001001: fsqrt_table = 23'b10000010111111010000011;
10'b0001001010: fsqrt_table = 23'b10000011010100011010101;
10'b0001001011: fsqrt_table = 23'b10000011101001100011101;
10'b0001001100: fsqrt_table = 23'b10000011111110101011100;
10'b0001001101: fsqrt_table = 23'b10000100010011110010010;
10'b0001001110: fsqrt_table = 23'b10000100101000110111111;
10'b0001001111: fsqrt_table = 23'b10000100111101111100011;
10'b0001010000: fsqrt_table = 23'b10000101010010111111110;
10'b0001010001: fsqrt_table = 23'b10000101101000000001111;
10'b0001010010: fsqrt_table = 23'b10000101111101000011000;
10'b0001010011: fsqrt_table = 23'b10000110010010000010111;
10'b0001010100: fsqrt_table = 23'b10000110100111000001101;
10'b0001010101: fsqrt_table = 23'b10000110111011111111011;
10'b0001010110: fsqrt_table = 23'b10000111010000111011111;
10'b0001010111: fsqrt_table = 23'b10000111100101110111010;
10'b0001011000: fsqrt_table = 23'b10000111111010110001101;
10'b0001011001: fsqrt_table = 23'b10001000001111101010110;
10'b0001011010: fsqrt_table = 23'b10001000100100100010111;
10'b0001011011: fsqrt_table = 23'b10001000111001011001111;
10'b0001011100: fsqrt_table = 23'b10001001001110001111110;
10'b0001011101: fsqrt_table = 23'b10001001100011000100100;
10'b0001011110: fsqrt_table = 23'b10001001110111111000001;
10'b0001011111: fsqrt_table = 23'b10001010001100101010101;
10'b0001100000: fsqrt_table = 23'b10001010100001011100001;
10'b0001100001: fsqrt_table = 23'b10001010110110001100100;
10'b0001100010: fsqrt_table = 23'b10001011001010111011110;
10'b0001100011: fsqrt_table = 23'b10001011011111101010000;
10'b0001100100: fsqrt_table = 23'b10001011110100010111001;
10'b0001100101: fsqrt_table = 23'b10001100001001000011001;
10'b0001100110: fsqrt_table = 23'b10001100011101101110001;
10'b0001100111: fsqrt_table = 23'b10001100110010011000000;
10'b0001101000: fsqrt_table = 23'b10001101000111000000110;
10'b0001101001: fsqrt_table = 23'b10001101011011101000100;
10'b0001101010: fsqrt_table = 23'b10001101110000001111001;
10'b0001101011: fsqrt_table = 23'b10001110000100110100110;
10'b0001101100: fsqrt_table = 23'b10001110011001011001010;
10'b0001101101: fsqrt_table = 23'b10001110101101111100110;
10'b0001101110: fsqrt_table = 23'b10001111000010011111001;
10'b0001101111: fsqrt_table = 23'b10001111010111000000100;
10'b0001110000: fsqrt_table = 23'b10001111101011100000110;
10'b0001110001: fsqrt_table = 23'b10010000000000000000000;
10'b0001110010: fsqrt_table = 23'b10010000010100011110010;
10'b0001110011: fsqrt_table = 23'b10010000101000111011011;
10'b0001110100: fsqrt_table = 23'b10010000111101010111100;
10'b0001110101: fsqrt_table = 23'b10010001010001110010100;
10'b0001110110: fsqrt_table = 23'b10010001100110001100100;
10'b0001110111: fsqrt_table = 23'b10010001111010100101100;
10'b0001111000: fsqrt_table = 23'b10010010001110111101100;
10'b0001111001: fsqrt_table = 23'b10010010100011010100011;
10'b0001111010: fsqrt_table = 23'b10010010110111101010011;
10'b0001111011: fsqrt_table = 23'b10010011001011111111001;
10'b0001111100: fsqrt_table = 23'b10010011100000010011000;
10'b0001111101: fsqrt_table = 23'b10010011110100100101111;
10'b0001111110: fsqrt_table = 23'b10010100001000110111101;
10'b0001111111: fsqrt_table = 23'b10010100011101001000100;
10'b0010000000: fsqrt_table = 23'b10010100110001011000010;
10'b0010000001: fsqrt_table = 23'b10010101000101100111000;
10'b0010000010: fsqrt_table = 23'b10010101011001110100110;
10'b0010000011: fsqrt_table = 23'b10010101101110000001100;
10'b0010000100: fsqrt_table = 23'b10010110000010001101010;
10'b0010000101: fsqrt_table = 23'b10010110010110011000000;
10'b0010000110: fsqrt_table = 23'b10010110101010100001110;
10'b0010000111: fsqrt_table = 23'b10010110111110101010100;
10'b0010001000: fsqrt_table = 23'b10010111010010110010010;
10'b0010001001: fsqrt_table = 23'b10010111100110111001000;
10'b0010001010: fsqrt_table = 23'b10010111111010111110110;
10'b0010001011: fsqrt_table = 23'b10011000001111000011100;
10'b0010001100: fsqrt_table = 23'b10011000100011000111010;
10'b0010001101: fsqrt_table = 23'b10011000110111001010001;
10'b0010001110: fsqrt_table = 23'b10011001001011001011111;
10'b0010001111: fsqrt_table = 23'b10011001011111001100110;
10'b0010010000: fsqrt_table = 23'b10011001110011001100101;
10'b0010010001: fsqrt_table = 23'b10011010000111001011100;
10'b0010010010: fsqrt_table = 23'b10011010011011001001011;
10'b0010010011: fsqrt_table = 23'b10011010101111000110011;
10'b0010010100: fsqrt_table = 23'b10011011000011000010011;
10'b0010010101: fsqrt_table = 23'b10011011010110111101011;
10'b0010010110: fsqrt_table = 23'b10011011101010110111011;
10'b0010010111: fsqrt_table = 23'b10011011111110110000100;
10'b0010011000: fsqrt_table = 23'b10011100010010101000101;
10'b0010011001: fsqrt_table = 23'b10011100100110011111110;
10'b0010011010: fsqrt_table = 23'b10011100111010010110000;
10'b0010011011: fsqrt_table = 23'b10011101001110001011010;
10'b0010011100: fsqrt_table = 23'b10011101100001111111100;
10'b0010011101: fsqrt_table = 23'b10011101110101110010111;
10'b0010011110: fsqrt_table = 23'b10011110001001100101010;
10'b0010011111: fsqrt_table = 23'b10011110011101010110110;
10'b0010100000: fsqrt_table = 23'b10011110110001000111010;
10'b0010100001: fsqrt_table = 23'b10011111000100110110111;
10'b0010100010: fsqrt_table = 23'b10011111011000100101100;
10'b0010100011: fsqrt_table = 23'b10011111101100010011010;
10'b0010100100: fsqrt_table = 23'b10100000000000000000000;
10'b0010100101: fsqrt_table = 23'b10100000010011101011111;
10'b0010100110: fsqrt_table = 23'b10100000100111010110110;
10'b0010100111: fsqrt_table = 23'b10100000111011000000110;
10'b0010101000: fsqrt_table = 23'b10100001001110101001110;
10'b0010101001: fsqrt_table = 23'b10100001100010010001111;
10'b0010101010: fsqrt_table = 23'b10100001110101111001001;
10'b0010101011: fsqrt_table = 23'b10100010001001011111011;
10'b0010101100: fsqrt_table = 23'b10100010011101000100110;
10'b0010101101: fsqrt_table = 23'b10100010110000101001010;
10'b0010101110: fsqrt_table = 23'b10100011000100001100110;
10'b0010101111: fsqrt_table = 23'b10100011010111101111100;
10'b0010110000: fsqrt_table = 23'b10100011101011010001001;
10'b0010110001: fsqrt_table = 23'b10100011111110110010000;
10'b0010110010: fsqrt_table = 23'b10100100010010010001111;
10'b0010110011: fsqrt_table = 23'b10100100100101110000111;
10'b0010110100: fsqrt_table = 23'b10100100111001001111000;
10'b0010110101: fsqrt_table = 23'b10100101001100101100010;
10'b0010110110: fsqrt_table = 23'b10100101100000001000100;
10'b0010110111: fsqrt_table = 23'b10100101110011100011111;
10'b0010111000: fsqrt_table = 23'b10100110000110111110011;
10'b0010111001: fsqrt_table = 23'b10100110011010011000000;
10'b0010111010: fsqrt_table = 23'b10100110101101110000110;
10'b0010111011: fsqrt_table = 23'b10100111000001001000101;
10'b0010111100: fsqrt_table = 23'b10100111010100011111101;
10'b0010111101: fsqrt_table = 23'b10100111100111110101101;
10'b0010111110: fsqrt_table = 23'b10100111111011001010111;
10'b0010111111: fsqrt_table = 23'b10101000001110011111001;
10'b0011000000: fsqrt_table = 23'b10101000100001110010101;
10'b0011000001: fsqrt_table = 23'b10101000110101000101001;
10'b0011000010: fsqrt_table = 23'b10101001001000010110110;
10'b0011000011: fsqrt_table = 23'b10101001011011100111101;
10'b0011000100: fsqrt_table = 23'b10101001101110110111100;
10'b0011000101: fsqrt_table = 23'b10101010000010000110101;
10'b0011000110: fsqrt_table = 23'b10101010010101010100110;
10'b0011000111: fsqrt_table = 23'b10101010101000100010001;
10'b0011001000: fsqrt_table = 23'b10101010111011101110101;
10'b0011001001: fsqrt_table = 23'b10101011001110111010010;
10'b0011001010: fsqrt_table = 23'b10101011100010000100111;
10'b0011001011: fsqrt_table = 23'b10101011110101001110111;
10'b0011001100: fsqrt_table = 23'b10101100001000010111111;
10'b0011001101: fsqrt_table = 23'b10101100011011100000000;
10'b0011001110: fsqrt_table = 23'b10101100101110100111011;
10'b0011001111: fsqrt_table = 23'b10101101000001101101110;
10'b0011010000: fsqrt_table = 23'b10101101010100110011011;
10'b0011010001: fsqrt_table = 23'b10101101100111111000001;
10'b0011010010: fsqrt_table = 23'b10101101111010111100001;
10'b0011010011: fsqrt_table = 23'b10101110001101111111001;
10'b0011010100: fsqrt_table = 23'b10101110100001000001011;
10'b0011010101: fsqrt_table = 23'b10101110110100000010110;
10'b0011010110: fsqrt_table = 23'b10101111000111000011011;
10'b0011010111: fsqrt_table = 23'b10101111011010000011001;
10'b0011011000: fsqrt_table = 23'b10101111101101000010000;
10'b0011011001: fsqrt_table = 23'b10110000000000000000000;
10'b0011011010: fsqrt_table = 23'b10110000010010111101010;
10'b0011011011: fsqrt_table = 23'b10110000100101111001101;
10'b0011011100: fsqrt_table = 23'b10110000111000110101001;
10'b0011011101: fsqrt_table = 23'b10110001001011101111111;
10'b0011011110: fsqrt_table = 23'b10110001011110101001110;
10'b0011011111: fsqrt_table = 23'b10110001110001100010111;
10'b0011100000: fsqrt_table = 23'b10110010000100011011001;
10'b0011100001: fsqrt_table = 23'b10110010010111010010100;
10'b0011100010: fsqrt_table = 23'b10110010101010001001001;
10'b0011100011: fsqrt_table = 23'b10110010111100111111000;
10'b0011100100: fsqrt_table = 23'b10110011001111110100000;
10'b0011100101: fsqrt_table = 23'b10110011100010101000001;
10'b0011100110: fsqrt_table = 23'b10110011110101011011100;
10'b0011100111: fsqrt_table = 23'b10110100001000001110000;
10'b0011101000: fsqrt_table = 23'b10110100011010111111110;
10'b0011101001: fsqrt_table = 23'b10110100101101110000101;
10'b0011101010: fsqrt_table = 23'b10110101000000100000110;
10'b0011101011: fsqrt_table = 23'b10110101010011010000001;
10'b0011101100: fsqrt_table = 23'b10110101100101111110101;
10'b0011101101: fsqrt_table = 23'b10110101111000101100011;
10'b0011101110: fsqrt_table = 23'b10110110001011011001010;
10'b0011101111: fsqrt_table = 23'b10110110011110000101011;
10'b0011110000: fsqrt_table = 23'b10110110110000110000110;
10'b0011110001: fsqrt_table = 23'b10110111000011011011010;
10'b0011110010: fsqrt_table = 23'b10110111010110000101000;
10'b0011110011: fsqrt_table = 23'b10110111101000101101111;
10'b0011110100: fsqrt_table = 23'b10110111111011010110001;
10'b0011110101: fsqrt_table = 23'b10111000001101111101100;
10'b0011110110: fsqrt_table = 23'b10111000100000100100000;
10'b0011110111: fsqrt_table = 23'b10111000110011001001111;
10'b0011111000: fsqrt_table = 23'b10111001000101101110111;
10'b0011111001: fsqrt_table = 23'b10111001011000010011001;
10'b0011111010: fsqrt_table = 23'b10111001101010110110100;
10'b0011111011: fsqrt_table = 23'b10111001111101011001001;
10'b0011111100: fsqrt_table = 23'b10111010001111111011001;
10'b0011111101: fsqrt_table = 23'b10111010100010011100010;
10'b0011111110: fsqrt_table = 23'b10111010110100111100100;
10'b0011111111: fsqrt_table = 23'b10111011000111011100001;
10'b0100000000: fsqrt_table = 23'b10111011011001111010111;
10'b0100000001: fsqrt_table = 23'b10111011101100011000111;
10'b0100000010: fsqrt_table = 23'b10111011111110110110010;
10'b0100000011: fsqrt_table = 23'b10111100010001010010110;
10'b0100000100: fsqrt_table = 23'b10111100100011101110011;
10'b0100000101: fsqrt_table = 23'b10111100110110001001011;
10'b0100000110: fsqrt_table = 23'b10111101001000100011101;
10'b0100000111: fsqrt_table = 23'b10111101011010111101000;
10'b0100001000: fsqrt_table = 23'b10111101101101010101110;
10'b0100001001: fsqrt_table = 23'b10111101111111101101101;
10'b0100001010: fsqrt_table = 23'b10111110010010000100110;
10'b0100001011: fsqrt_table = 23'b10111110100100011011010;
10'b0100001100: fsqrt_table = 23'b10111110110110110000111;
10'b0100001101: fsqrt_table = 23'b10111111001001000101110;
10'b0100001110: fsqrt_table = 23'b10111111011011011001111;
10'b0100001111: fsqrt_table = 23'b10111111101101101101011;
10'b0100010000: fsqrt_table = 23'b11000000000000000000000;
10'b0100010001: fsqrt_table = 23'b11000000010010010001111;
10'b0100010010: fsqrt_table = 23'b11000000100100100011001;
10'b0100010011: fsqrt_table = 23'b11000000110110110011100;
10'b0100010100: fsqrt_table = 23'b11000001001001000011001;
10'b0100010101: fsqrt_table = 23'b11000001011011010010001;
10'b0100010110: fsqrt_table = 23'b11000001101101100000011;
10'b0100010111: fsqrt_table = 23'b11000001111111101101110;
10'b0100011000: fsqrt_table = 23'b11000010010001111010100;
10'b0100011001: fsqrt_table = 23'b11000010100100000110100;
10'b0100011010: fsqrt_table = 23'b11000010110110010001110;
10'b0100011011: fsqrt_table = 23'b11000011001000011100010;
10'b0100011100: fsqrt_table = 23'b11000011011010100110001;
10'b0100011101: fsqrt_table = 23'b11000011101100101111001;
10'b0100011110: fsqrt_table = 23'b11000011111110110111100;
10'b0100011111: fsqrt_table = 23'b11000100010000111111001;
10'b0100100000: fsqrt_table = 23'b11000100100011000110000;
10'b0100100001: fsqrt_table = 23'b11000100110101001100001;
10'b0100100010: fsqrt_table = 23'b11000101000111010001101;
10'b0100100011: fsqrt_table = 23'b11000101011001010110011;
10'b0100100100: fsqrt_table = 23'b11000101101011011010011;
10'b0100100101: fsqrt_table = 23'b11000101111101011101101;
10'b0100100110: fsqrt_table = 23'b11000110001111100000001;
10'b0100100111: fsqrt_table = 23'b11000110100001100010000;
10'b0100101000: fsqrt_table = 23'b11000110110011100011001;
10'b0100101001: fsqrt_table = 23'b11000111000101100011100;
10'b0100101010: fsqrt_table = 23'b11000111010111100011010;
10'b0100101011: fsqrt_table = 23'b11000111101001100010010;
10'b0100101100: fsqrt_table = 23'b11000111111011100000100;
10'b0100101101: fsqrt_table = 23'b11001000001101011110001;
10'b0100101110: fsqrt_table = 23'b11001000011111011011000;
10'b0100101111: fsqrt_table = 23'b11001000110001010111001;
10'b0100110000: fsqrt_table = 23'b11001001000011010010101;
10'b0100110001: fsqrt_table = 23'b11001001010101001101011;
10'b0100110010: fsqrt_table = 23'b11001001100111000111011;
10'b0100110011: fsqrt_table = 23'b11001001111001000000110;
10'b0100110100: fsqrt_table = 23'b11001010001010111001100;
10'b0100110101: fsqrt_table = 23'b11001010011100110001011;
10'b0100110110: fsqrt_table = 23'b11001010101110101000101;
10'b0100110111: fsqrt_table = 23'b11001011000000011111010;
10'b0100111000: fsqrt_table = 23'b11001011010010010101001;
10'b0100111001: fsqrt_table = 23'b11001011100100001010010;
10'b0100111010: fsqrt_table = 23'b11001011110101111110110;
10'b0100111011: fsqrt_table = 23'b11001100000111110010101;
10'b0100111100: fsqrt_table = 23'b11001100011001100101110;
10'b0100111101: fsqrt_table = 23'b11001100101011011000001;
10'b0100111110: fsqrt_table = 23'b11001100111101001001111;
10'b0100111111: fsqrt_table = 23'b11001101001110111010111;
10'b0101000000: fsqrt_table = 23'b11001101100000101011010;
10'b0101000001: fsqrt_table = 23'b11001101110010011011000;
10'b0101000010: fsqrt_table = 23'b11001110000100001010000;
10'b0101000011: fsqrt_table = 23'b11001110010101111000010;
10'b0101000100: fsqrt_table = 23'b11001110100111100101111;
10'b0101000101: fsqrt_table = 23'b11001110111001010010111;
10'b0101000110: fsqrt_table = 23'b11001111001010111111001;
10'b0101000111: fsqrt_table = 23'b11001111011100101010110;
10'b0101001000: fsqrt_table = 23'b11001111101110010101110;
10'b0101001001: fsqrt_table = 23'b11010000000000000000000;
10'b0101001010: fsqrt_table = 23'b11010000010001101001101;
10'b0101001011: fsqrt_table = 23'b11010000100011010010100;
10'b0101001100: fsqrt_table = 23'b11010000110100111010110;
10'b0101001101: fsqrt_table = 23'b11010001000110100010011;
10'b0101001110: fsqrt_table = 23'b11010001011000001001010;
10'b0101001111: fsqrt_table = 23'b11010001101001101111100;
10'b0101010000: fsqrt_table = 23'b11010001111011010101001;
10'b0101010001: fsqrt_table = 23'b11010010001100111010000;
10'b0101010010: fsqrt_table = 23'b11010010011110011110011;
10'b0101010011: fsqrt_table = 23'b11010010110000000001111;
10'b0101010100: fsqrt_table = 23'b11010011000001100100111;
10'b0101010101: fsqrt_table = 23'b11010011010011000111001;
10'b0101010110: fsqrt_table = 23'b11010011100100101000110;
10'b0101010111: fsqrt_table = 23'b11010011110110001001110;
10'b0101011000: fsqrt_table = 23'b11010100000111101010000;
10'b0101011001: fsqrt_table = 23'b11010100011001001001110;
10'b0101011010: fsqrt_table = 23'b11010100101010101000110;
10'b0101011011: fsqrt_table = 23'b11010100111100000111001;
10'b0101011100: fsqrt_table = 23'b11010101001101100100110;
10'b0101011101: fsqrt_table = 23'b11010101011111000001111;
10'b0101011110: fsqrt_table = 23'b11010101110000011110010;
10'b0101011111: fsqrt_table = 23'b11010110000001111010000;
10'b0101100000: fsqrt_table = 23'b11010110010011010101001;
10'b0101100001: fsqrt_table = 23'b11010110100100101111101;
10'b0101100010: fsqrt_table = 23'b11010110110110001001011;
10'b0101100011: fsqrt_table = 23'b11010111000111100010101;
10'b0101100100: fsqrt_table = 23'b11010111011000111011001;
10'b0101100101: fsqrt_table = 23'b11010111101010010011000;
10'b0101100110: fsqrt_table = 23'b11010111111011101010010;
10'b0101100111: fsqrt_table = 23'b11011000001101000000111;
10'b0101101000: fsqrt_table = 23'b11011000011110010110111;
10'b0101101001: fsqrt_table = 23'b11011000101111101100010;
10'b0101101010: fsqrt_table = 23'b11011001000001000001000;
10'b0101101011: fsqrt_table = 23'b11011001010010010101000;
10'b0101101100: fsqrt_table = 23'b11011001100011101000100;
10'b0101101101: fsqrt_table = 23'b11011001110100111011010;
10'b0101101110: fsqrt_table = 23'b11011010000110001101100;
10'b0101101111: fsqrt_table = 23'b11011010010111011111000;
10'b0101110000: fsqrt_table = 23'b11011010101000101111111;
10'b0101110001: fsqrt_table = 23'b11011010111010000000010;
10'b0101110010: fsqrt_table = 23'b11011011001011001111111;
10'b0101110011: fsqrt_table = 23'b11011011011100011111000;
10'b0101110100: fsqrt_table = 23'b11011011101101101101011;
10'b0101110101: fsqrt_table = 23'b11011011111110111011001;
10'b0101110110: fsqrt_table = 23'b11011100010000001000011;
10'b0101110111: fsqrt_table = 23'b11011100100001010100111;
10'b0101111000: fsqrt_table = 23'b11011100110010100000111;
10'b0101111001: fsqrt_table = 23'b11011101000011101100001;
10'b0101111010: fsqrt_table = 23'b11011101010100110110111;
10'b0101111011: fsqrt_table = 23'b11011101100110000000111;
10'b0101111100: fsqrt_table = 23'b11011101110111001010011;
10'b0101111101: fsqrt_table = 23'b11011110001000010011010;
10'b0101111110: fsqrt_table = 23'b11011110011001011011100;
10'b0101111111: fsqrt_table = 23'b11011110101010100011000;
10'b0110000000: fsqrt_table = 23'b11011110111011101010001;
10'b0110000001: fsqrt_table = 23'b11011111001100110000100;
10'b0110000010: fsqrt_table = 23'b11011111011101110110010;
10'b0110000011: fsqrt_table = 23'b11011111101110111011011;
10'b0110000100: fsqrt_table = 23'b11100000000000000000000;
10'b0110000101: fsqrt_table = 23'b11100000010001000100000;
10'b0110000110: fsqrt_table = 23'b11100000100010000111011;
10'b0110000111: fsqrt_table = 23'b11100000110011001010001;
10'b0110001000: fsqrt_table = 23'b11100001000100001100010;
10'b0110001001: fsqrt_table = 23'b11100001010101001101110;
10'b0110001010: fsqrt_table = 23'b11100001100110001110110;
10'b0110001011: fsqrt_table = 23'b11100001110111001111000;
10'b0110001100: fsqrt_table = 23'b11100010001000001110110;
10'b0110001101: fsqrt_table = 23'b11100010011001001110000;
10'b0110001110: fsqrt_table = 23'b11100010101010001100100;
10'b0110001111: fsqrt_table = 23'b11100010111011001010100;
10'b0110010000: fsqrt_table = 23'b11100011001100000111110;
10'b0110010001: fsqrt_table = 23'b11100011011101000100100;
10'b0110010010: fsqrt_table = 23'b11100011101110000000110;
10'b0110010011: fsqrt_table = 23'b11100011111110111100010;
10'b0110010100: fsqrt_table = 23'b11100100001111110111010;
10'b0110010101: fsqrt_table = 23'b11100100100000110001101;
10'b0110010110: fsqrt_table = 23'b11100100110001101011100;
10'b0110010111: fsqrt_table = 23'b11100101000010100100101;
10'b0110011000: fsqrt_table = 23'b11100101010011011101010;
10'b0110011001: fsqrt_table = 23'b11100101100100010101011;
10'b0110011010: fsqrt_table = 23'b11100101110101001100110;
10'b0110011011: fsqrt_table = 23'b11100110000110000011101;
10'b0110011100: fsqrt_table = 23'b11100110010110111001111;
10'b0110011101: fsqrt_table = 23'b11100110100111101111101;
10'b0110011110: fsqrt_table = 23'b11100110111000100100110;
10'b0110011111: fsqrt_table = 23'b11100111001001011001010;
10'b0110100000: fsqrt_table = 23'b11100111011010001101010;
10'b0110100001: fsqrt_table = 23'b11100111101011000000101;
10'b0110100010: fsqrt_table = 23'b11100111111011110011011;
10'b0110100011: fsqrt_table = 23'b11101000001100100101101;
10'b0110100100: fsqrt_table = 23'b11101000011101010111010;
10'b0110100101: fsqrt_table = 23'b11101000101110001000010;
10'b0110100110: fsqrt_table = 23'b11101000111110111000110;
10'b0110100111: fsqrt_table = 23'b11101001001111101000110;
10'b0110101000: fsqrt_table = 23'b11101001100000011000000;
10'b0110101001: fsqrt_table = 23'b11101001110001000110111;
10'b0110101010: fsqrt_table = 23'b11101010000001110101000;
10'b0110101011: fsqrt_table = 23'b11101010010010100010101;
10'b0110101100: fsqrt_table = 23'b11101010100011001111110;
10'b0110101101: fsqrt_table = 23'b11101010110011111100010;
10'b0110101110: fsqrt_table = 23'b11101011000100101000001;
10'b0110101111: fsqrt_table = 23'b11101011010101010011100;
10'b0110110000: fsqrt_table = 23'b11101011100101111110010;
10'b0110110001: fsqrt_table = 23'b11101011110110101000100;
10'b0110110010: fsqrt_table = 23'b11101100000111010010001;
10'b0110110011: fsqrt_table = 23'b11101100010111111011010;
10'b0110110100: fsqrt_table = 23'b11101100101000100011110;
10'b0110110101: fsqrt_table = 23'b11101100111001001011110;
10'b0110110110: fsqrt_table = 23'b11101101001001110011001;
10'b0110110111: fsqrt_table = 23'b11101101011010011010000;
10'b0110111000: fsqrt_table = 23'b11101101101011000000011;
10'b0110111001: fsqrt_table = 23'b11101101111011100110001;
10'b0110111010: fsqrt_table = 23'b11101110001100001011010;
10'b0110111011: fsqrt_table = 23'b11101110011100101111111;
10'b0110111100: fsqrt_table = 23'b11101110101101010100000;
10'b0110111101: fsqrt_table = 23'b11101110111101110111100;
10'b0110111110: fsqrt_table = 23'b11101111001110011010011;
10'b0110111111: fsqrt_table = 23'b11101111011110111100111;
10'b0111000000: fsqrt_table = 23'b11101111101111011110110;
10'b0111000001: fsqrt_table = 23'b11110000000000000000000;
10'b0111000010: fsqrt_table = 23'b11110000010000100000110;
10'b0111000011: fsqrt_table = 23'b11110000100001000001000;
10'b0111000100: fsqrt_table = 23'b11110000110001100000101;
10'b0111000101: fsqrt_table = 23'b11110001000001111111110;
10'b0111000110: fsqrt_table = 23'b11110001010010011110010;
10'b0111000111: fsqrt_table = 23'b11110001100010111100011;
10'b0111001000: fsqrt_table = 23'b11110001110011011001110;
10'b0111001001: fsqrt_table = 23'b11110010000011110110110;
10'b0111001010: fsqrt_table = 23'b11110010010100010011001;
10'b0111001011: fsqrt_table = 23'b11110010100100101111000;
10'b0111001100: fsqrt_table = 23'b11110010110101001010010;
10'b0111001101: fsqrt_table = 23'b11110011000101100101000;
10'b0111001110: fsqrt_table = 23'b11110011010101111111010;
10'b0111001111: fsqrt_table = 23'b11110011100110011001000;
10'b0111010000: fsqrt_table = 23'b11110011110110110010001;
10'b0111010001: fsqrt_table = 23'b11110100000111001010110;
10'b0111010010: fsqrt_table = 23'b11110100010111100010110;
10'b0111010011: fsqrt_table = 23'b11110100100111111010010;
10'b0111010100: fsqrt_table = 23'b11110100111000010001011;
10'b0111010101: fsqrt_table = 23'b11110101001000100111110;
10'b0111010110: fsqrt_table = 23'b11110101011000111101110;
10'b0111010111: fsqrt_table = 23'b11110101101001010011001;
10'b0111011000: fsqrt_table = 23'b11110101111001101000000;
10'b0111011001: fsqrt_table = 23'b11110110001001111100011;
10'b0111011010: fsqrt_table = 23'b11110110011010010000001;
10'b0111011011: fsqrt_table = 23'b11110110101010100011011;
10'b0111011100: fsqrt_table = 23'b11110110111010110110001;
10'b0111011101: fsqrt_table = 23'b11110111001011001000011;
10'b0111011110: fsqrt_table = 23'b11110111011011011010001;
10'b0111011111: fsqrt_table = 23'b11110111101011101011010;
10'b0111100000: fsqrt_table = 23'b11110111111011111011111;
10'b0111100001: fsqrt_table = 23'b11111000001100001100000;
10'b0111100010: fsqrt_table = 23'b11111000011100011011101;
10'b0111100011: fsqrt_table = 23'b11111000101100101010110;
10'b0111100100: fsqrt_table = 23'b11111000111100111001010;
10'b0111100101: fsqrt_table = 23'b11111001001101000111010;
10'b0111100110: fsqrt_table = 23'b11111001011101010100111;
10'b0111100111: fsqrt_table = 23'b11111001101101100001111;
10'b0111101000: fsqrt_table = 23'b11111001111101101110010;
10'b0111101001: fsqrt_table = 23'b11111010001101111010010;
10'b0111101010: fsqrt_table = 23'b11111010011110000101101;
10'b0111101011: fsqrt_table = 23'b11111010101110010000101;
10'b0111101100: fsqrt_table = 23'b11111010111110011011000;
10'b0111101101: fsqrt_table = 23'b11111011001110100100111;
10'b0111101110: fsqrt_table = 23'b11111011011110101110010;
10'b0111101111: fsqrt_table = 23'b11111011101110110111001;
10'b0111110000: fsqrt_table = 23'b11111011111110111111100;
10'b0111110001: fsqrt_table = 23'b11111100001111000111011;
10'b0111110010: fsqrt_table = 23'b11111100011111001110101;
10'b0111110011: fsqrt_table = 23'b11111100101111010101100;
10'b0111110100: fsqrt_table = 23'b11111100111111011011110;
10'b0111110101: fsqrt_table = 23'b11111101001111100001101;
10'b0111110110: fsqrt_table = 23'b11111101011111100110111;
10'b0111110111: fsqrt_table = 23'b11111101101111101011101;
10'b0111111000: fsqrt_table = 23'b11111101111111101111111;
10'b0111111001: fsqrt_table = 23'b11111110001111110011110;
10'b0111111010: fsqrt_table = 23'b11111110011111110111000;
10'b0111111011: fsqrt_table = 23'b11111110101111111001110;
10'b0111111100: fsqrt_table = 23'b11111110111111111100000;
10'b0111111101: fsqrt_table = 23'b11111111001111111101110;
10'b0111111110: fsqrt_table = 23'b11111111011111111111000;
10'b0111111111: fsqrt_table = 23'b11111111101111111111110;
10'b1000000000: fsqrt_table = 23'b00000000000000000000000;
10'b1000000001: fsqrt_table = 23'b00000000001111111111100;
10'b1000000010: fsqrt_table = 23'b00000000011111111110000;
10'b1000000011: fsqrt_table = 23'b00000000101111111011100;
10'b1000000100: fsqrt_table = 23'b00000000111111111000000;
10'b1000000101: fsqrt_table = 23'b00000001001111110011100;
10'b1000000110: fsqrt_table = 23'b00000001011111101110001;
10'b1000000111: fsqrt_table = 23'b00000001101111100111101;
10'b1000001000: fsqrt_table = 23'b00000001111111100000010;
10'b1000001001: fsqrt_table = 23'b00000010001111010111111;
10'b1000001010: fsqrt_table = 23'b00000010011111001110100;
10'b1000001011: fsqrt_table = 23'b00000010101111000100001;
10'b1000001100: fsqrt_table = 23'b00000010111110111000111;
10'b1000001101: fsqrt_table = 23'b00000011001110101100100;
10'b1000001110: fsqrt_table = 23'b00000011011110011111011;
10'b1000001111: fsqrt_table = 23'b00000011101110010001001;
10'b1000010000: fsqrt_table = 23'b00000011111110000010000;
10'b1000010001: fsqrt_table = 23'b00000100001101110001111;
10'b1000010010: fsqrt_table = 23'b00000100011101100000110;
10'b1000010011: fsqrt_table = 23'b00000100101101001110110;
10'b1000010100: fsqrt_table = 23'b00000100111100111011111;
10'b1000010101: fsqrt_table = 23'b00000101001100100111111;
10'b1000010110: fsqrt_table = 23'b00000101011100010011001;
10'b1000010111: fsqrt_table = 23'b00000101101011111101010;
10'b1000011000: fsqrt_table = 23'b00000101111011100110100;
10'b1000011001: fsqrt_table = 23'b00000110001011001110111;
10'b1000011010: fsqrt_table = 23'b00000110011010110110011;
10'b1000011011: fsqrt_table = 23'b00000110101010011100110;
10'b1000011100: fsqrt_table = 23'b00000110111010000010011;
10'b1000011101: fsqrt_table = 23'b00000111001001100111000;
10'b1000011110: fsqrt_table = 23'b00000111011001001010110;
10'b1000011111: fsqrt_table = 23'b00000111101000101101100;
10'b1000100000: fsqrt_table = 23'b00000111111000001111011;
10'b1000100001: fsqrt_table = 23'b00001000000111110000011;
10'b1000100010: fsqrt_table = 23'b00001000010111010000011;
10'b1000100011: fsqrt_table = 23'b00001000100110101111101;
10'b1000100100: fsqrt_table = 23'b00001000110110001101111;
10'b1000100101: fsqrt_table = 23'b00001001000101101011001;
10'b1000100110: fsqrt_table = 23'b00001001010101000111101;
10'b1000100111: fsqrt_table = 23'b00001001100100100011001;
10'b1000101000: fsqrt_table = 23'b00001001110011111101110;
10'b1000101001: fsqrt_table = 23'b00001010000011010111100;
10'b1000101010: fsqrt_table = 23'b00001010010010110000011;
10'b1000101011: fsqrt_table = 23'b00001010100010001000011;
10'b1000101100: fsqrt_table = 23'b00001010110001011111100;
10'b1000101101: fsqrt_table = 23'b00001011000000110101110;
10'b1000101110: fsqrt_table = 23'b00001011010000001011000;
10'b1000101111: fsqrt_table = 23'b00001011011111011111100;
10'b1000110000: fsqrt_table = 23'b00001011101110110011000;
10'b1000110001: fsqrt_table = 23'b00001011111110000101110;
10'b1000110010: fsqrt_table = 23'b00001100001101010111100;
10'b1000110011: fsqrt_table = 23'b00001100011100101000100;
10'b1000110100: fsqrt_table = 23'b00001100101011111000101;
10'b1000110101: fsqrt_table = 23'b00001100111011000111110;
10'b1000110110: fsqrt_table = 23'b00001101001010010110001;
10'b1000110111: fsqrt_table = 23'b00001101011001100011101;
10'b1000111000: fsqrt_table = 23'b00001101101000110000010;
10'b1000111001: fsqrt_table = 23'b00001101110111111100001;
10'b1000111010: fsqrt_table = 23'b00001110000111000111000;
10'b1000111011: fsqrt_table = 23'b00001110010110010001001;
10'b1000111100: fsqrt_table = 23'b00001110100101011010011;
10'b1000111101: fsqrt_table = 23'b00001110110100100010110;
10'b1000111110: fsqrt_table = 23'b00001111000011101010010;
10'b1000111111: fsqrt_table = 23'b00001111010010110001000;
10'b1001000000: fsqrt_table = 23'b00001111100001110110110;
10'b1001000001: fsqrt_table = 23'b00001111110000111011111;
10'b1001000010: fsqrt_table = 23'b00010000000000000000000;
10'b1001000011: fsqrt_table = 23'b00010000001111000011011;
10'b1001000100: fsqrt_table = 23'b00010000011110000101111;
10'b1001000101: fsqrt_table = 23'b00010000101101000111100;
10'b1001000110: fsqrt_table = 23'b00010000111100001000011;
10'b1001000111: fsqrt_table = 23'b00010001001011001000100;
10'b1001001000: fsqrt_table = 23'b00010001011010000111101;
10'b1001001001: fsqrt_table = 23'b00010001101001000110000;
10'b1001001010: fsqrt_table = 23'b00010001111000000011101;
10'b1001001011: fsqrt_table = 23'b00010010000111000000011;
10'b1001001100: fsqrt_table = 23'b00010010010101111100011;
10'b1001001101: fsqrt_table = 23'b00010010100100110111100;
10'b1001001110: fsqrt_table = 23'b00010010110011110001110;
10'b1001001111: fsqrt_table = 23'b00010011000010101011010;
10'b1001010000: fsqrt_table = 23'b00010011010001100100000;
10'b1001010001: fsqrt_table = 23'b00010011100000011011111;
10'b1001010010: fsqrt_table = 23'b00010011101111010011000;
10'b1001010011: fsqrt_table = 23'b00010011111110001001010;
10'b1001010100: fsqrt_table = 23'b00010100001100111110110;
10'b1001010101: fsqrt_table = 23'b00010100011011110011100;
10'b1001010110: fsqrt_table = 23'b00010100101010100111011;
10'b1001010111: fsqrt_table = 23'b00010100111001011010100;
10'b1001011000: fsqrt_table = 23'b00010101001000001100111;
10'b1001011001: fsqrt_table = 23'b00010101010110111110011;
10'b1001011010: fsqrt_table = 23'b00010101100101101111001;
10'b1001011011: fsqrt_table = 23'b00010101110100011111001;
10'b1001011100: fsqrt_table = 23'b00010110000011001110010;
10'b1001011101: fsqrt_table = 23'b00010110010001111100101;
10'b1001011110: fsqrt_table = 23'b00010110100000101010010;
10'b1001011111: fsqrt_table = 23'b00010110101111010111001;
10'b1001100000: fsqrt_table = 23'b00010110111110000011010;
10'b1001100001: fsqrt_table = 23'b00010111001100101110100;
10'b1001100010: fsqrt_table = 23'b00010111011011011001000;
10'b1001100011: fsqrt_table = 23'b00010111101010000010110;
10'b1001100100: fsqrt_table = 23'b00010111111000101011110;
10'b1001100101: fsqrt_table = 23'b00011000000111010100000;
10'b1001100110: fsqrt_table = 23'b00011000010101111011100;
10'b1001100111: fsqrt_table = 23'b00011000100100100010010;
10'b1001101000: fsqrt_table = 23'b00011000110011001000001;
10'b1001101001: fsqrt_table = 23'b00011001000001101101011;
10'b1001101010: fsqrt_table = 23'b00011001010000010001110;
10'b1001101011: fsqrt_table = 23'b00011001011110110101011;
10'b1001101100: fsqrt_table = 23'b00011001101101011000011;
10'b1001101101: fsqrt_table = 23'b00011001111011111010100;
10'b1001101110: fsqrt_table = 23'b00011010001010011100000;
10'b1001101111: fsqrt_table = 23'b00011010011000111100101;
10'b1001110000: fsqrt_table = 23'b00011010100111011100100;
10'b1001110001: fsqrt_table = 23'b00011010110101111011110;
10'b1001110010: fsqrt_table = 23'b00011011000100011010010;
10'b1001110011: fsqrt_table = 23'b00011011010010110111111;
10'b1001110100: fsqrt_table = 23'b00011011100001010100111;
10'b1001110101: fsqrt_table = 23'b00011011101111110001001;
10'b1001110110: fsqrt_table = 23'b00011011111110001100101;
10'b1001110111: fsqrt_table = 23'b00011100001100100111011;
10'b1001111000: fsqrt_table = 23'b00011100011011000001011;
10'b1001111001: fsqrt_table = 23'b00011100101001011010110;
10'b1001111010: fsqrt_table = 23'b00011100110111110011010;
10'b1001111011: fsqrt_table = 23'b00011101000110001011001;
10'b1001111100: fsqrt_table = 23'b00011101010100100010010;
10'b1001111101: fsqrt_table = 23'b00011101100010111000110;
10'b1001111110: fsqrt_table = 23'b00011101110001001110011;
10'b1001111111: fsqrt_table = 23'b00011101111111100011011;
10'b1010000000: fsqrt_table = 23'b00011110001101110111101;
10'b1010000001: fsqrt_table = 23'b00011110011100001011001;
10'b1010000010: fsqrt_table = 23'b00011110101010011110000;
10'b1010000011: fsqrt_table = 23'b00011110111000110000001;
10'b1010000100: fsqrt_table = 23'b00011111000111000001100;
10'b1010000101: fsqrt_table = 23'b00011111010101010010001;
10'b1010000110: fsqrt_table = 23'b00011111100011100010001;
10'b1010000111: fsqrt_table = 23'b00011111110001110001011;
10'b1010001000: fsqrt_table = 23'b00100000000000000000000;
10'b1010001001: fsqrt_table = 23'b00100000001110001101111;
10'b1010001010: fsqrt_table = 23'b00100000011100011011000;
10'b1010001011: fsqrt_table = 23'b00100000101010100111100;
10'b1010001100: fsqrt_table = 23'b00100000111000110011010;
10'b1010001101: fsqrt_table = 23'b00100001000110111110011;
10'b1010001110: fsqrt_table = 23'b00100001010101001000110;
10'b1010001111: fsqrt_table = 23'b00100001100011010010100;
10'b1010010000: fsqrt_table = 23'b00100001110001011011100;
10'b1010010001: fsqrt_table = 23'b00100001111111100011110;
10'b1010010010: fsqrt_table = 23'b00100010001101101011011;
10'b1010010011: fsqrt_table = 23'b00100010011011110010010;
10'b1010010100: fsqrt_table = 23'b00100010101001111000100;
10'b1010010101: fsqrt_table = 23'b00100010110111111110001;
10'b1010010110: fsqrt_table = 23'b00100011000110000011000;
10'b1010010111: fsqrt_table = 23'b00100011010100000111010;
10'b1010011000: fsqrt_table = 23'b00100011100010001010110;
10'b1010011001: fsqrt_table = 23'b00100011110000001101101;
10'b1010011010: fsqrt_table = 23'b00100011111110001111110;
10'b1010011011: fsqrt_table = 23'b00100100001100010001010;
10'b1010011100: fsqrt_table = 23'b00100100011010010010001;
10'b1010011101: fsqrt_table = 23'b00100100101000010010010;
10'b1010011110: fsqrt_table = 23'b00100100110110010001110;
10'b1010011111: fsqrt_table = 23'b00100101000100010000101;
10'b1010100000: fsqrt_table = 23'b00100101010010001110110;
10'b1010100001: fsqrt_table = 23'b00100101100000001100010;
10'b1010100010: fsqrt_table = 23'b00100101101110001001000;
10'b1010100011: fsqrt_table = 23'b00100101111100000101010;
10'b1010100100: fsqrt_table = 23'b00100110001010000000110;
10'b1010100101: fsqrt_table = 23'b00100110010111111011100;
10'b1010100110: fsqrt_table = 23'b00100110100101110101110;
10'b1010100111: fsqrt_table = 23'b00100110110011101111010;
10'b1010101000: fsqrt_table = 23'b00100111000001101000001;
10'b1010101001: fsqrt_table = 23'b00100111001111100000011;
10'b1010101010: fsqrt_table = 23'b00100111011101010111111;
10'b1010101011: fsqrt_table = 23'b00100111101011001110111;
10'b1010101100: fsqrt_table = 23'b00100111111001000101001;
10'b1010101101: fsqrt_table = 23'b00101000000110111010110;
10'b1010101110: fsqrt_table = 23'b00101000010100101111110;
10'b1010101111: fsqrt_table = 23'b00101000100010100100000;
10'b1010110000: fsqrt_table = 23'b00101000110000010111110;
10'b1010110001: fsqrt_table = 23'b00101000111110001010110;
10'b1010110010: fsqrt_table = 23'b00101001001011111101001;
10'b1010110011: fsqrt_table = 23'b00101001011001101111000;
10'b1010110100: fsqrt_table = 23'b00101001100111100000001;
10'b1010110101: fsqrt_table = 23'b00101001110101010000100;
10'b1010110110: fsqrt_table = 23'b00101010000011000000011;
10'b1010110111: fsqrt_table = 23'b00101010010000101111101;
10'b1010111000: fsqrt_table = 23'b00101010011110011110010;
10'b1010111001: fsqrt_table = 23'b00101010101100001100001;
10'b1010111010: fsqrt_table = 23'b00101010111001111001100;
10'b1010111011: fsqrt_table = 23'b00101011000111100110010;
10'b1010111100: fsqrt_table = 23'b00101011010101010010010;
10'b1010111101: fsqrt_table = 23'b00101011100010111101110;
10'b1010111110: fsqrt_table = 23'b00101011110000101000101;
10'b1010111111: fsqrt_table = 23'b00101011111110010010110;
10'b1011000000: fsqrt_table = 23'b00101100001011111100011;
10'b1011000001: fsqrt_table = 23'b00101100011001100101010;
10'b1011000010: fsqrt_table = 23'b00101100100111001101101;
10'b1011000011: fsqrt_table = 23'b00101100110100110101011;
10'b1011000100: fsqrt_table = 23'b00101101000010011100100;
10'b1011000101: fsqrt_table = 23'b00101101010000000011000;
10'b1011000110: fsqrt_table = 23'b00101101011101101000111;
10'b1011000111: fsqrt_table = 23'b00101101101011001110001;
10'b1011001000: fsqrt_table = 23'b00101101111000110010110;
10'b1011001001: fsqrt_table = 23'b00101110000110010110111;
10'b1011001010: fsqrt_table = 23'b00101110010011111010010;
10'b1011001011: fsqrt_table = 23'b00101110100001011101001;
10'b1011001100: fsqrt_table = 23'b00101110101110111111010;
10'b1011001101: fsqrt_table = 23'b00101110111100100000111;
10'b1011001110: fsqrt_table = 23'b00101111001010000010000;
10'b1011001111: fsqrt_table = 23'b00101111010111100010011;
10'b1011010000: fsqrt_table = 23'b00101111100101000010001;
10'b1011010001: fsqrt_table = 23'b00101111110010100001011;
10'b1011010010: fsqrt_table = 23'b00110000000000000000000;
10'b1011010011: fsqrt_table = 23'b00110000001101011110000;
10'b1011010100: fsqrt_table = 23'b00110000011010111011100;
10'b1011010101: fsqrt_table = 23'b00110000101000011000010;
10'b1011010110: fsqrt_table = 23'b00110000110101110100100;
10'b1011010111: fsqrt_table = 23'b00110001000011010000001;
10'b1011011000: fsqrt_table = 23'b00110001010000101011010;
10'b1011011001: fsqrt_table = 23'b00110001011110000101101;
10'b1011011010: fsqrt_table = 23'b00110001101011011111100;
10'b1011011011: fsqrt_table = 23'b00110001111000111000110;
10'b1011011100: fsqrt_table = 23'b00110010000110010001100;
10'b1011011101: fsqrt_table = 23'b00110010010011101001101;
10'b1011011110: fsqrt_table = 23'b00110010100001000001001;
10'b1011011111: fsqrt_table = 23'b00110010101110011000001;
10'b1011100000: fsqrt_table = 23'b00110010111011101110100;
10'b1011100001: fsqrt_table = 23'b00110011001001000100010;
10'b1011100010: fsqrt_table = 23'b00110011010110011001100;
10'b1011100011: fsqrt_table = 23'b00110011100011101110001;
10'b1011100100: fsqrt_table = 23'b00110011110001000010001;
10'b1011100101: fsqrt_table = 23'b00110011111110010101101;
10'b1011100110: fsqrt_table = 23'b00110100001011101000100;
10'b1011100111: fsqrt_table = 23'b00110100011000111010111;
10'b1011101000: fsqrt_table = 23'b00110100100110001100101;
10'b1011101001: fsqrt_table = 23'b00110100110011011101110;
10'b1011101010: fsqrt_table = 23'b00110101000000101110011;
10'b1011101011: fsqrt_table = 23'b00110101001101111110100;
10'b1011101100: fsqrt_table = 23'b00110101011011001101111;
10'b1011101101: fsqrt_table = 23'b00110101101000011100111;
10'b1011101110: fsqrt_table = 23'b00110101110101101011001;
10'b1011101111: fsqrt_table = 23'b00110110000010111001000;
10'b1011110000: fsqrt_table = 23'b00110110010000000110010;
10'b1011110001: fsqrt_table = 23'b00110110011101010010111;
10'b1011110010: fsqrt_table = 23'b00110110101010011111000;
10'b1011110011: fsqrt_table = 23'b00110110110111101010100;
10'b1011110100: fsqrt_table = 23'b00110111000100110101100;
10'b1011110101: fsqrt_table = 23'b00110111010001111111111;
10'b1011110110: fsqrt_table = 23'b00110111011111001001110;
10'b1011110111: fsqrt_table = 23'b00110111101100010011001;
10'b1011111000: fsqrt_table = 23'b00110111111001011011111;
10'b1011111001: fsqrt_table = 23'b00111000000110100100000;
10'b1011111010: fsqrt_table = 23'b00111000010011101011101;
10'b1011111011: fsqrt_table = 23'b00111000100000110010110;
10'b1011111100: fsqrt_table = 23'b00111000101101111001011;
10'b1011111101: fsqrt_table = 23'b00111000111010111111011;
10'b1011111110: fsqrt_table = 23'b00111001001000000100110;
10'b1011111111: fsqrt_table = 23'b00111001010101001001110;
10'b1100000000: fsqrt_table = 23'b00111001100010001110001;
10'b1100000001: fsqrt_table = 23'b00111001101111010001111;
10'b1100000010: fsqrt_table = 23'b00111001111100010101001;
10'b1100000011: fsqrt_table = 23'b00111010001001010111111;
10'b1100000100: fsqrt_table = 23'b00111010010110011010001;
10'b1100000101: fsqrt_table = 23'b00111010100011011011110;
10'b1100000110: fsqrt_table = 23'b00111010110000011100111;
10'b1100000111: fsqrt_table = 23'b00111010111101011101100;
10'b1100001000: fsqrt_table = 23'b00111011001010011101100;
10'b1100001001: fsqrt_table = 23'b00111011010111011101000;
10'b1100001010: fsqrt_table = 23'b00111011100100011100000;
10'b1100001011: fsqrt_table = 23'b00111011110001011010011;
10'b1100001100: fsqrt_table = 23'b00111011111110011000010;
10'b1100001101: fsqrt_table = 23'b00111100001011010101101;
10'b1100001110: fsqrt_table = 23'b00111100011000010010100;
10'b1100001111: fsqrt_table = 23'b00111100100101001110111;
10'b1100010000: fsqrt_table = 23'b00111100110010001010101;
10'b1100010001: fsqrt_table = 23'b00111100111111000101111;
10'b1100010010: fsqrt_table = 23'b00111101001100000000101;
10'b1100010011: fsqrt_table = 23'b00111101011000111010110;
10'b1100010100: fsqrt_table = 23'b00111101100101110100100;
10'b1100010101: fsqrt_table = 23'b00111101110010101101101;
10'b1100010110: fsqrt_table = 23'b00111101111111100110010;
10'b1100010111: fsqrt_table = 23'b00111110001100011110011;
10'b1100011000: fsqrt_table = 23'b00111110011001010101111;
10'b1100011001: fsqrt_table = 23'b00111110100110001101000;
10'b1100011010: fsqrt_table = 23'b00111110110011000011100;
10'b1100011011: fsqrt_table = 23'b00111110111111111001101;
10'b1100011100: fsqrt_table = 23'b00111111001100101111001;
10'b1100011101: fsqrt_table = 23'b00111111011001100100001;
10'b1100011110: fsqrt_table = 23'b00111111100110011000101;
10'b1100011111: fsqrt_table = 23'b00111111110011001100100;
10'b1100100000: fsqrt_table = 23'b01000000000000000000000;
10'b1100100001: fsqrt_table = 23'b01000000001100110011000;
10'b1100100010: fsqrt_table = 23'b01000000011001100101011;
10'b1100100011: fsqrt_table = 23'b01000000100110010111010;
10'b1100100100: fsqrt_table = 23'b01000000110011001000110;
10'b1100100101: fsqrt_table = 23'b01000000111111111001101;
10'b1100100110: fsqrt_table = 23'b01000001001100101010000;
10'b1100100111: fsqrt_table = 23'b01000001011001011001111;
10'b1100101000: fsqrt_table = 23'b01000001100110001001010;
10'b1100101001: fsqrt_table = 23'b01000001110010111000001;
10'b1100101010: fsqrt_table = 23'b01000001111111100110100;
10'b1100101011: fsqrt_table = 23'b01000010001100010100011;
10'b1100101100: fsqrt_table = 23'b01000010011001000001110;
10'b1100101101: fsqrt_table = 23'b01000010100101101110101;
10'b1100101110: fsqrt_table = 23'b01000010110010011011000;
10'b1100101111: fsqrt_table = 23'b01000010111111000110111;
10'b1100110000: fsqrt_table = 23'b01000011001011110010010;
10'b1100110001: fsqrt_table = 23'b01000011011000011101010;
10'b1100110010: fsqrt_table = 23'b01000011100101000111101;
10'b1100110011: fsqrt_table = 23'b01000011110001110001100;
10'b1100110100: fsqrt_table = 23'b01000011111110011010111;
10'b1100110101: fsqrt_table = 23'b01000100001011000011110;
10'b1100110110: fsqrt_table = 23'b01000100010111101100001;
10'b1100110111: fsqrt_table = 23'b01000100100100010100001;
10'b1100111000: fsqrt_table = 23'b01000100110000111011100;
10'b1100111001: fsqrt_table = 23'b01000100111101100010100;
10'b1100111010: fsqrt_table = 23'b01000101001010001000111;
10'b1100111011: fsqrt_table = 23'b01000101010110101110111;
10'b1100111100: fsqrt_table = 23'b01000101100011010100011;
10'b1100111101: fsqrt_table = 23'b01000101101111111001011;
10'b1100111110: fsqrt_table = 23'b01000101111100011101111;
10'b1100111111: fsqrt_table = 23'b01000110001001000001111;
10'b1101000000: fsqrt_table = 23'b01000110010101100101011;
10'b1101000001: fsqrt_table = 23'b01000110100010001000011;
10'b1101000010: fsqrt_table = 23'b01000110101110101011000;
10'b1101000011: fsqrt_table = 23'b01000110111011001101001;
10'b1101000100: fsqrt_table = 23'b01000111000111101110101;
10'b1101000101: fsqrt_table = 23'b01000111010100001111111;
10'b1101000110: fsqrt_table = 23'b01000111100000110000100;
10'b1101000111: fsqrt_table = 23'b01000111101101010000101;
10'b1101001000: fsqrt_table = 23'b01000111111001110000011;
10'b1101001001: fsqrt_table = 23'b01001000000110001111100;
10'b1101001010: fsqrt_table = 23'b01001000010010101110010;
10'b1101001011: fsqrt_table = 23'b01001000011111001100101;
10'b1101001100: fsqrt_table = 23'b01001000101011101010011;
10'b1101001101: fsqrt_table = 23'b01001000111000000111101;
10'b1101001110: fsqrt_table = 23'b01001001000100100100100;
10'b1101001111: fsqrt_table = 23'b01001001010001000000111;
10'b1101010000: fsqrt_table = 23'b01001001011101011100111;
10'b1101010001: fsqrt_table = 23'b01001001101001111000010;
10'b1101010010: fsqrt_table = 23'b01001001110110010011010;
10'b1101010011: fsqrt_table = 23'b01001010000010101101110;
10'b1101010100: fsqrt_table = 23'b01001010001111000111110;
10'b1101010101: fsqrt_table = 23'b01001010011011100001011;
10'b1101010110: fsqrt_table = 23'b01001010100111111010100;
10'b1101010111: fsqrt_table = 23'b01001010110100010011001;
10'b1101011000: fsqrt_table = 23'b01001011000000101011010;
10'b1101011001: fsqrt_table = 23'b01001011001101000011000;
10'b1101011010: fsqrt_table = 23'b01001011011001011010010;
10'b1101011011: fsqrt_table = 23'b01001011100101110001001;
10'b1101011100: fsqrt_table = 23'b01001011110010000111011;
10'b1101011101: fsqrt_table = 23'b01001011111110011101010;
10'b1101011110: fsqrt_table = 23'b01001100001010110010110;
10'b1101011111: fsqrt_table = 23'b01001100010111000111101;
10'b1101100000: fsqrt_table = 23'b01001100100011011100001;
10'b1101100001: fsqrt_table = 23'b01001100101111110000010;
10'b1101100010: fsqrt_table = 23'b01001100111100000011111;
10'b1101100011: fsqrt_table = 23'b01001101001000010111000;
10'b1101100100: fsqrt_table = 23'b01001101010100101001101;
10'b1101100101: fsqrt_table = 23'b01001101100000111011111;
10'b1101100110: fsqrt_table = 23'b01001101101101001101101;
10'b1101100111: fsqrt_table = 23'b01001101111001011111000;
10'b1101101000: fsqrt_table = 23'b01001110000101101111111;
10'b1101101001: fsqrt_table = 23'b01001110010010000000010;
10'b1101101010: fsqrt_table = 23'b01001110011110010000010;
10'b1101101011: fsqrt_table = 23'b01001110101010011111110;
10'b1101101100: fsqrt_table = 23'b01001110110110101110111;
10'b1101101101: fsqrt_table = 23'b01001111000010111101100;
10'b1101101110: fsqrt_table = 23'b01001111001111001011110;
10'b1101101111: fsqrt_table = 23'b01001111011011011001011;
10'b1101110000: fsqrt_table = 23'b01001111100111100110110;
10'b1101110001: fsqrt_table = 23'b01001111110011110011101;
10'b1101110010: fsqrt_table = 23'b01010000000000000000000;
10'b1101110011: fsqrt_table = 23'b01010000001100001100000;
10'b1101110100: fsqrt_table = 23'b01010000011000010111100;
10'b1101110101: fsqrt_table = 23'b01010000100100100010101;
10'b1101110110: fsqrt_table = 23'b01010000110000101101010;
10'b1101110111: fsqrt_table = 23'b01010000111100110111100;
10'b1101111000: fsqrt_table = 23'b01010001001001000001010;
10'b1101111001: fsqrt_table = 23'b01010001010101001010100;
10'b1101111010: fsqrt_table = 23'b01010001100001010011011;
10'b1101111011: fsqrt_table = 23'b01010001101101011011111;
10'b1101111100: fsqrt_table = 23'b01010001111001100011111;
10'b1101111101: fsqrt_table = 23'b01010010000101101011100;
10'b1101111110: fsqrt_table = 23'b01010010010001110010101;
10'b1101111111: fsqrt_table = 23'b01010010011101111001011;
10'b1110000000: fsqrt_table = 23'b01010010101001111111101;
10'b1110000001: fsqrt_table = 23'b01010010110110000101100;
10'b1110000010: fsqrt_table = 23'b01010011000010001011000;
10'b1110000011: fsqrt_table = 23'b01010011001110001111111;
10'b1110000100: fsqrt_table = 23'b01010011011010010100100;
10'b1110000101: fsqrt_table = 23'b01010011100110011000101;
10'b1110000110: fsqrt_table = 23'b01010011110010011100011;
10'b1110000111: fsqrt_table = 23'b01010011111110011111101;
10'b1110001000: fsqrt_table = 23'b01010100001010100010100;
10'b1110001001: fsqrt_table = 23'b01010100010110100100111;
10'b1110001010: fsqrt_table = 23'b01010100100010100110111;
10'b1110001011: fsqrt_table = 23'b01010100101110101000100;
10'b1110001100: fsqrt_table = 23'b01010100111010101001101;
10'b1110001101: fsqrt_table = 23'b01010101000110101010011;
10'b1110001110: fsqrt_table = 23'b01010101010010101010101;
10'b1110001111: fsqrt_table = 23'b01010101011110101010100;
10'b1110010000: fsqrt_table = 23'b01010101101010101010000;
10'b1110010001: fsqrt_table = 23'b01010101110110101001000;
10'b1110010010: fsqrt_table = 23'b01010110000010100111101;
10'b1110010011: fsqrt_table = 23'b01010110001110100101111;
10'b1110010100: fsqrt_table = 23'b01010110011010100011101;
10'b1110010101: fsqrt_table = 23'b01010110100110100001000;
10'b1110010110: fsqrt_table = 23'b01010110110010011110000;
10'b1110010111: fsqrt_table = 23'b01010110111110011010100;
10'b1110011000: fsqrt_table = 23'b01010111001010010110101;
10'b1110011001: fsqrt_table = 23'b01010111010110010010010;
10'b1110011010: fsqrt_table = 23'b01010111100010001101101;
10'b1110011011: fsqrt_table = 23'b01010111101110001000100;
10'b1110011100: fsqrt_table = 23'b01010111111010000010111;
10'b1110011101: fsqrt_table = 23'b01011000000101111101000;
10'b1110011110: fsqrt_table = 23'b01011000010001110110101;
10'b1110011111: fsqrt_table = 23'b01011000011101101111111;
10'b1110100000: fsqrt_table = 23'b01011000101001101000101;
10'b1110100001: fsqrt_table = 23'b01011000110101100001000;
10'b1110100010: fsqrt_table = 23'b01011001000001011001000;
10'b1110100011: fsqrt_table = 23'b01011001001101010000101;
10'b1110100100: fsqrt_table = 23'b01011001011001000111110;
10'b1110100101: fsqrt_table = 23'b01011001100100111110101;
10'b1110100110: fsqrt_table = 23'b01011001110000110101000;
10'b1110100111: fsqrt_table = 23'b01011001111100101010111;
10'b1110101000: fsqrt_table = 23'b01011010001000100000100;
10'b1110101001: fsqrt_table = 23'b01011010010100010101101;
10'b1110101010: fsqrt_table = 23'b01011010100000001010011;
10'b1110101011: fsqrt_table = 23'b01011010101011111110101;
10'b1110101100: fsqrt_table = 23'b01011010110111110010101;
10'b1110101101: fsqrt_table = 23'b01011011000011100110001;
10'b1110101110: fsqrt_table = 23'b01011011001111011001010;
10'b1110101111: fsqrt_table = 23'b01011011011011001100000;
10'b1110110000: fsqrt_table = 23'b01011011100110111110011;
10'b1110110001: fsqrt_table = 23'b01011011110010110000010;
10'b1110110010: fsqrt_table = 23'b01011011111110100001111;
10'b1110110011: fsqrt_table = 23'b01011100001010010011000;
10'b1110110100: fsqrt_table = 23'b01011100010110000011110;
10'b1110110101: fsqrt_table = 23'b01011100100001110100000;
10'b1110110110: fsqrt_table = 23'b01011100101101100100000;
10'b1110110111: fsqrt_table = 23'b01011100111001010011100;
10'b1110111000: fsqrt_table = 23'b01011101000101000010110;
10'b1110111001: fsqrt_table = 23'b01011101010000110001100;
10'b1110111010: fsqrt_table = 23'b01011101011100011111111;
10'b1110111011: fsqrt_table = 23'b01011101101000001101111;
10'b1110111100: fsqrt_table = 23'b01011101110011111011011;
10'b1110111101: fsqrt_table = 23'b01011101111111101000101;
10'b1110111110: fsqrt_table = 23'b01011110001011010101011;
10'b1110111111: fsqrt_table = 23'b01011110010111000001110;
10'b1111000000: fsqrt_table = 23'b01011110100010101101111;
10'b1111000001: fsqrt_table = 23'b01011110101110011001100;
10'b1111000010: fsqrt_table = 23'b01011110111010000100110;
10'b1111000011: fsqrt_table = 23'b01011111000101101111100;
10'b1111000100: fsqrt_table = 23'b01011111010001011010000;
10'b1111000101: fsqrt_table = 23'b01011111011101000100001;
10'b1111000110: fsqrt_table = 23'b01011111101000101101110;
10'b1111000111: fsqrt_table = 23'b01011111110100010111001;
10'b1111001000: fsqrt_table = 23'b01100000000000000000000;
10'b1111001001: fsqrt_table = 23'b01100000001011101000100;
10'b1111001010: fsqrt_table = 23'b01100000010111010000101;
10'b1111001011: fsqrt_table = 23'b01100000100010111000100;
10'b1111001100: fsqrt_table = 23'b01100000101110011111111;
10'b1111001101: fsqrt_table = 23'b01100000111010000110111;
10'b1111001110: fsqrt_table = 23'b01100001000101101101100;
10'b1111001111: fsqrt_table = 23'b01100001010001010011110;
10'b1111010000: fsqrt_table = 23'b01100001011100111001100;
10'b1111010001: fsqrt_table = 23'b01100001101000011111000;
10'b1111010010: fsqrt_table = 23'b01100001110100000100001;
10'b1111010011: fsqrt_table = 23'b01100001111111101000111;
10'b1111010100: fsqrt_table = 23'b01100010001011001101010;
10'b1111010101: fsqrt_table = 23'b01100010010110110001001;
10'b1111010110: fsqrt_table = 23'b01100010100010010100110;
10'b1111010111: fsqrt_table = 23'b01100010101101111000000;
10'b1111011000: fsqrt_table = 23'b01100010111001011010110;
10'b1111011001: fsqrt_table = 23'b01100011000100111101010;
10'b1111011010: fsqrt_table = 23'b01100011010000011111011;
10'b1111011011: fsqrt_table = 23'b01100011011100000001000;
10'b1111011100: fsqrt_table = 23'b01100011100111100010011;
10'b1111011101: fsqrt_table = 23'b01100011110011000011011;
10'b1111011110: fsqrt_table = 23'b01100011111110100100000;
10'b1111011111: fsqrt_table = 23'b01100100001010000100001;
10'b1111100000: fsqrt_table = 23'b01100100010101100100000;
10'b1111100001: fsqrt_table = 23'b01100100100001000011100;
10'b1111100010: fsqrt_table = 23'b01100100101100100010101;
10'b1111100011: fsqrt_table = 23'b01100100111000000001011;
10'b1111100100: fsqrt_table = 23'b01100101000011011111110;
10'b1111100101: fsqrt_table = 23'b01100101001110111101110;
10'b1111100110: fsqrt_table = 23'b01100101011010011011011;
10'b1111100111: fsqrt_table = 23'b01100101100101111000101;
10'b1111101000: fsqrt_table = 23'b01100101110001010101100;
10'b1111101001: fsqrt_table = 23'b01100101111100110010000;
10'b1111101010: fsqrt_table = 23'b01100110001000001110010;
10'b1111101011: fsqrt_table = 23'b01100110010011101010000;
10'b1111101100: fsqrt_table = 23'b01100110011111000101100;
10'b1111101101: fsqrt_table = 23'b01100110101010100000100;
10'b1111101110: fsqrt_table = 23'b01100110110101111011010;
10'b1111101111: fsqrt_table = 23'b01100111000001010101101;
10'b1111110000: fsqrt_table = 23'b01100111001100101111100;
10'b1111110001: fsqrt_table = 23'b01100111011000001001001;
10'b1111110010: fsqrt_table = 23'b01100111100011100010011;
10'b1111110011: fsqrt_table = 23'b01100111101110111011011;
10'b1111110100: fsqrt_table = 23'b01100111111010010011111;
10'b1111110101: fsqrt_table = 23'b01101000000101101100000;
10'b1111110110: fsqrt_table = 23'b01101000010001000011111;
10'b1111110111: fsqrt_table = 23'b01101000011100011011011;
10'b1111111000: fsqrt_table = 23'b01101000100111110010011;
10'b1111111001: fsqrt_table = 23'b01101000110011001001001;
10'b1111111010: fsqrt_table = 23'b01101000111110011111100;
10'b1111111011: fsqrt_table = 23'b01101001001001110101101;
10'b1111111100: fsqrt_table = 23'b01101001010101001011010;
10'b1111111101: fsqrt_table = 23'b01101001100000100000101;
10'b1111111110: fsqrt_table = 23'b01101001101011110101100;
10'b1111111111: fsqrt_table = 23'b01101001110111001010001;

     endcase
    end
  endfunction

  function [22:0] fsqrtinv_table (
    input [9:0] e_m2 );
    begin
      case(e_m2)

10'b0000000000: fsqrtinv_table = 23'b01101010000010011110011;
10'b0000000001: fsqrtinv_table = 23'b01101001101011111000011;
10'b0000000010: fsqrtinv_table = 23'b01101001010101010110100;
10'b0000000011: fsqrtinv_table = 23'b01101000111110111000111;
10'b0000000100: fsqrtinv_table = 23'b01101000101000011111100;
10'b0000000101: fsqrtinv_table = 23'b01101000010010001010010;
10'b0000000110: fsqrtinv_table = 23'b01100111111011111001001;
10'b0000000111: fsqrtinv_table = 23'b01100111100101101100001;
10'b0000001000: fsqrtinv_table = 23'b01100111001111100011001;
10'b0000001001: fsqrtinv_table = 23'b01100110111001011110011;
10'b0000001010: fsqrtinv_table = 23'b01100110100011011101101;
10'b0000001011: fsqrtinv_table = 23'b01100110001101100000111;
10'b0000001100: fsqrtinv_table = 23'b01100101110111101000001;
10'b0000001101: fsqrtinv_table = 23'b01100101100001110011100;
10'b0000001110: fsqrtinv_table = 23'b01100101001100000010110;
10'b0000001111: fsqrtinv_table = 23'b01100100110110010110000;
10'b0000010000: fsqrtinv_table = 23'b01100100100000101101010;
10'b0000010001: fsqrtinv_table = 23'b01100100001011001000011;
10'b0000010010: fsqrtinv_table = 23'b01100011110101100111011;
10'b0000010011: fsqrtinv_table = 23'b01100011100000001010011;
10'b0000010100: fsqrtinv_table = 23'b01100011001010110001001;
10'b0000010101: fsqrtinv_table = 23'b01100010110101011011110;
10'b0000010110: fsqrtinv_table = 23'b01100010100000001010010;
10'b0000010111: fsqrtinv_table = 23'b01100010001010111100101;
10'b0000011000: fsqrtinv_table = 23'b01100001110101110010110;
10'b0000011001: fsqrtinv_table = 23'b01100001100000101100101;
10'b0000011010: fsqrtinv_table = 23'b01100001001011101010010;
10'b0000011011: fsqrtinv_table = 23'b01100000110110101011110;
10'b0000011100: fsqrtinv_table = 23'b01100000100001110000111;
10'b0000011101: fsqrtinv_table = 23'b01100000001100111001110;
10'b0000011110: fsqrtinv_table = 23'b01011111111000000110010;
10'b0000011111: fsqrtinv_table = 23'b01011111100011010110100;
10'b0000100000: fsqrtinv_table = 23'b01011111001110101010011;
10'b0000100001: fsqrtinv_table = 23'b01011110111010000010000;
10'b0000100010: fsqrtinv_table = 23'b01011110100101011101001;
10'b0000100011: fsqrtinv_table = 23'b01011110010000111011111;
10'b0000100100: fsqrtinv_table = 23'b01011101111100011110010;
10'b0000100101: fsqrtinv_table = 23'b01011101101000000100010;
10'b0000100110: fsqrtinv_table = 23'b01011101010011101101110;
10'b0000100111: fsqrtinv_table = 23'b01011100111111011010111;
10'b0000101000: fsqrtinv_table = 23'b01011100101011001011100;
10'b0000101001: fsqrtinv_table = 23'b01011100010110111111101;
10'b0000101010: fsqrtinv_table = 23'b01011100000010110111010;
10'b0000101011: fsqrtinv_table = 23'b01011011101110110010011;
10'b0000101100: fsqrtinv_table = 23'b01011011011010110000111;
10'b0000101101: fsqrtinv_table = 23'b01011011000110110010111;
10'b0000101110: fsqrtinv_table = 23'b01011010110010111000011;
10'b0000101111: fsqrtinv_table = 23'b01011010011111000001010;
10'b0000110000: fsqrtinv_table = 23'b01011010001011001101100;
10'b0000110001: fsqrtinv_table = 23'b01011001110111011101010;
10'b0000110010: fsqrtinv_table = 23'b01011001100011110000010;
10'b0000110011: fsqrtinv_table = 23'b01011001010000000110110;
10'b0000110100: fsqrtinv_table = 23'b01011000111100100000100;
10'b0000110101: fsqrtinv_table = 23'b01011000101000111101101;
10'b0000110110: fsqrtinv_table = 23'b01011000010101011110000;
10'b0000110111: fsqrtinv_table = 23'b01011000000010000001110;
10'b0000111000: fsqrtinv_table = 23'b01010111101110101000110;
10'b0000111001: fsqrtinv_table = 23'b01010111011011010011000;
10'b0000111010: fsqrtinv_table = 23'b01010111001000000000100;
10'b0000111011: fsqrtinv_table = 23'b01010110110100110001010;
10'b0000111100: fsqrtinv_table = 23'b01010110100001100101010;
10'b0000111101: fsqrtinv_table = 23'b01010110001110011100100;
10'b0000111110: fsqrtinv_table = 23'b01010101111011010110111;
10'b0000111111: fsqrtinv_table = 23'b01010101101000010100100;
10'b0001000000: fsqrtinv_table = 23'b01010101010101010101011;
10'b0001000001: fsqrtinv_table = 23'b01010101000010011001010;
10'b0001000010: fsqrtinv_table = 23'b01010100101111100000011;
10'b0001000011: fsqrtinv_table = 23'b01010100011100101010101;
10'b0001000100: fsqrtinv_table = 23'b01010100001001111000000;
10'b0001000101: fsqrtinv_table = 23'b01010011110111001000011;
10'b0001000110: fsqrtinv_table = 23'b01010011100100011100000;
10'b0001000111: fsqrtinv_table = 23'b01010011010001110010101;
10'b0001001000: fsqrtinv_table = 23'b01010010111111001100010;
10'b0001001001: fsqrtinv_table = 23'b01010010101100101001000;
10'b0001001010: fsqrtinv_table = 23'b01010010011010001000110;
10'b0001001011: fsqrtinv_table = 23'b01010010000111101011101;
10'b0001001100: fsqrtinv_table = 23'b01010001110101010001100;
10'b0001001101: fsqrtinv_table = 23'b01010001100010111010010;
10'b0001001110: fsqrtinv_table = 23'b01010001010000100110001;
10'b0001001111: fsqrtinv_table = 23'b01010000111110010100111;
10'b0001010000: fsqrtinv_table = 23'b01010000101100000110101;
10'b0001010001: fsqrtinv_table = 23'b01010000011001111011011;
10'b0001010010: fsqrtinv_table = 23'b01010000000111110011000;
10'b0001010011: fsqrtinv_table = 23'b01001111110101101101101;
10'b0001010100: fsqrtinv_table = 23'b01001111100011101011001;
10'b0001010101: fsqrtinv_table = 23'b01001111010001101011100;
10'b0001010110: fsqrtinv_table = 23'b01001110111111101110110;
10'b0001010111: fsqrtinv_table = 23'b01001110101101110100111;
10'b0001011000: fsqrtinv_table = 23'b01001110011011111110000;
10'b0001011001: fsqrtinv_table = 23'b01001110001010001001111;
10'b0001011010: fsqrtinv_table = 23'b01001101111000011000100;
10'b0001011011: fsqrtinv_table = 23'b01001101100110101010001;
10'b0001011100: fsqrtinv_table = 23'b01001101010100111110100;
10'b0001011101: fsqrtinv_table = 23'b01001101000011010101101;
10'b0001011110: fsqrtinv_table = 23'b01001100110001101111101;
10'b0001011111: fsqrtinv_table = 23'b01001100100000001100011;
10'b0001100000: fsqrtinv_table = 23'b01001100001110101011111;
10'b0001100001: fsqrtinv_table = 23'b01001011111101001110010;
10'b0001100010: fsqrtinv_table = 23'b01001011101011110011010;
10'b0001100011: fsqrtinv_table = 23'b01001011011010011011000;
10'b0001100100: fsqrtinv_table = 23'b01001011001001000101100;
10'b0001100101: fsqrtinv_table = 23'b01001010110111110010110;
10'b0001100110: fsqrtinv_table = 23'b01001010100110100010101;
10'b0001100111: fsqrtinv_table = 23'b01001010010101010101010;
10'b0001101000: fsqrtinv_table = 23'b01001010000100001010101;
10'b0001101001: fsqrtinv_table = 23'b01001001110011000010101;
10'b0001101010: fsqrtinv_table = 23'b01001001100001111101010;
10'b0001101011: fsqrtinv_table = 23'b01001001010000111010100;
10'b0001101100: fsqrtinv_table = 23'b01001000111111111010011;
10'b0001101101: fsqrtinv_table = 23'b01001000101110111101000;
10'b0001101110: fsqrtinv_table = 23'b01001000011110000010001;
10'b0001101111: fsqrtinv_table = 23'b01001000001101001001111;
10'b0001110000: fsqrtinv_table = 23'b01000111111100010100010;
10'b0001110001: fsqrtinv_table = 23'b01000111101011100001010;
10'b0001110010: fsqrtinv_table = 23'b01000111011010110000111;
10'b0001110011: fsqrtinv_table = 23'b01000111001010000010111;
10'b0001110100: fsqrtinv_table = 23'b01000110111001010111101;
10'b0001110101: fsqrtinv_table = 23'b01000110101000101110111;
10'b0001110110: fsqrtinv_table = 23'b01000110011000001000101;
10'b0001110111: fsqrtinv_table = 23'b01000110000111100100111;
10'b0001111000: fsqrtinv_table = 23'b01000101110111000011101;
10'b0001111001: fsqrtinv_table = 23'b01000101100110100101000;
10'b0001111010: fsqrtinv_table = 23'b01000101010110001000110;
10'b0001111011: fsqrtinv_table = 23'b01000101000101101111000;
10'b0001111100: fsqrtinv_table = 23'b01000100110101010111110;
10'b0001111101: fsqrtinv_table = 23'b01000100100101000011000;
10'b0001111110: fsqrtinv_table = 23'b01000100010100110000101;
10'b0001111111: fsqrtinv_table = 23'b01000100000100100000111;
10'b0010000000: fsqrtinv_table = 23'b01000011110100010011011;
10'b0010000001: fsqrtinv_table = 23'b01000011100100001000011;
10'b0010000010: fsqrtinv_table = 23'b01000011010011111111110;
10'b0010000011: fsqrtinv_table = 23'b01000011000011111001101;
10'b0010000100: fsqrtinv_table = 23'b01000010110011110101111;
10'b0010000101: fsqrtinv_table = 23'b01000010100011110100100;
10'b0010000110: fsqrtinv_table = 23'b01000010010011110101100;
10'b0010000111: fsqrtinv_table = 23'b01000010000011111000111;
10'b0010001000: fsqrtinv_table = 23'b01000001110011111110101;
10'b0010001001: fsqrtinv_table = 23'b01000001100100000110101;
10'b0010001010: fsqrtinv_table = 23'b01000001010100010001001;
10'b0010001011: fsqrtinv_table = 23'b01000001000100011101111;
10'b0010001100: fsqrtinv_table = 23'b01000000110100101101000;
10'b0010001101: fsqrtinv_table = 23'b01000000100100111110011;
10'b0010001110: fsqrtinv_table = 23'b01000000010101010010001;
10'b0010001111: fsqrtinv_table = 23'b01000000000101101000001;
10'b0010010000: fsqrtinv_table = 23'b00111111110110000000100;
10'b0010010001: fsqrtinv_table = 23'b00111111100110011011001;
10'b0010010010: fsqrtinv_table = 23'b00111111010110111000000;
10'b0010010011: fsqrtinv_table = 23'b00111111000111010111001;
10'b0010010100: fsqrtinv_table = 23'b00111110110111111000100;
10'b0010010101: fsqrtinv_table = 23'b00111110101000011100001;
10'b0010010110: fsqrtinv_table = 23'b00111110011001000010000;
10'b0010010111: fsqrtinv_table = 23'b00111110001001101010001;
10'b0010011000: fsqrtinv_table = 23'b00111101111010010100100;
10'b0010011001: fsqrtinv_table = 23'b00111101101011000001000;
10'b0010011010: fsqrtinv_table = 23'b00111101011011101111111;
10'b0010011011: fsqrtinv_table = 23'b00111101001100100000110;
10'b0010011100: fsqrtinv_table = 23'b00111100111101010100000;
10'b0010011101: fsqrtinv_table = 23'b00111100101110001001010;
10'b0010011110: fsqrtinv_table = 23'b00111100011111000000110;
10'b0010011111: fsqrtinv_table = 23'b00111100001111111010100;
10'b0010100000: fsqrtinv_table = 23'b00111100000000110110011;
10'b0010100001: fsqrtinv_table = 23'b00111011110001110100010;
10'b0010100010: fsqrtinv_table = 23'b00111011100010110100011;
10'b0010100011: fsqrtinv_table = 23'b00111011010011110110110;
10'b0010100100: fsqrtinv_table = 23'b00111011000100111011001;
10'b0010100101: fsqrtinv_table = 23'b00111010110110000001101;
10'b0010100110: fsqrtinv_table = 23'b00111010100111001010010;
10'b0010100111: fsqrtinv_table = 23'b00111010011000010100111;
10'b0010101000: fsqrtinv_table = 23'b00111010001001100001110;
10'b0010101001: fsqrtinv_table = 23'b00111001111010110000101;
10'b0010101010: fsqrtinv_table = 23'b00111001101100000001101;
10'b0010101011: fsqrtinv_table = 23'b00111001011101010100101;
10'b0010101100: fsqrtinv_table = 23'b00111001001110101001110;
10'b0010101101: fsqrtinv_table = 23'b00111001000000000001000;
10'b0010101110: fsqrtinv_table = 23'b00111000110001011010001;
10'b0010101111: fsqrtinv_table = 23'b00111000100010110101011;
10'b0010110000: fsqrtinv_table = 23'b00111000010100010010110;
10'b0010110001: fsqrtinv_table = 23'b00111000000101110010000;
10'b0010110010: fsqrtinv_table = 23'b00110111110111010011011;
10'b0010110011: fsqrtinv_table = 23'b00110111101000110110110;
10'b0010110100: fsqrtinv_table = 23'b00110111011010011100001;
10'b0010110101: fsqrtinv_table = 23'b00110111001100000011100;
10'b0010110110: fsqrtinv_table = 23'b00110110111101101100111;
10'b0010110111: fsqrtinv_table = 23'b00110110101111011000001;
10'b0010111000: fsqrtinv_table = 23'b00110110100001000101100;
10'b0010111001: fsqrtinv_table = 23'b00110110010010110100110;
10'b0010111010: fsqrtinv_table = 23'b00110110000100100110000;
10'b0010111011: fsqrtinv_table = 23'b00110101110110011001001;
10'b0010111100: fsqrtinv_table = 23'b00110101101000001110011;
10'b0010111101: fsqrtinv_table = 23'b00110101011010000101011;
10'b0010111110: fsqrtinv_table = 23'b00110101001011111110011;
10'b0010111111: fsqrtinv_table = 23'b00110100111101111001011;
10'b0011000000: fsqrtinv_table = 23'b00110100101111110110010;
10'b0011000001: fsqrtinv_table = 23'b00110100100001110101000;
10'b0011000010: fsqrtinv_table = 23'b00110100010011110101110;
10'b0011000011: fsqrtinv_table = 23'b00110100000101111000010;
10'b0011000100: fsqrtinv_table = 23'b00110011110111111100110;
10'b0011000101: fsqrtinv_table = 23'b00110011101010000011001;
10'b0011000110: fsqrtinv_table = 23'b00110011011100001011011;
10'b0011000111: fsqrtinv_table = 23'b00110011001110010101100;
10'b0011001000: fsqrtinv_table = 23'b00110011000000100001100;
10'b0011001001: fsqrtinv_table = 23'b00110010110010101111011;
10'b0011001010: fsqrtinv_table = 23'b00110010100100111111000;
10'b0011001011: fsqrtinv_table = 23'b00110010010111010000101;
10'b0011001100: fsqrtinv_table = 23'b00110010001001100100000;
10'b0011001101: fsqrtinv_table = 23'b00110001111011111001010;
10'b0011001110: fsqrtinv_table = 23'b00110001101110010000010;
10'b0011001111: fsqrtinv_table = 23'b00110001100000101001001;
10'b0011010000: fsqrtinv_table = 23'b00110001010011000011111;
10'b0011010001: fsqrtinv_table = 23'b00110001000101100000011;
10'b0011010010: fsqrtinv_table = 23'b00110000110111111110101;
10'b0011010011: fsqrtinv_table = 23'b00110000101010011110110;
10'b0011010100: fsqrtinv_table = 23'b00110000011101000000101;
10'b0011010101: fsqrtinv_table = 23'b00110000001111100100011;
10'b0011010110: fsqrtinv_table = 23'b00110000000010001001110;
10'b0011010111: fsqrtinv_table = 23'b00101111110100110001000;
10'b0011011000: fsqrtinv_table = 23'b00101111100111011010000;
10'b0011011001: fsqrtinv_table = 23'b00101111011010000100110;
10'b0011011010: fsqrtinv_table = 23'b00101111001100110001010;
10'b0011011011: fsqrtinv_table = 23'b00101110111111011111100;
10'b0011011100: fsqrtinv_table = 23'b00101110110010001111100;
10'b0011011101: fsqrtinv_table = 23'b00101110100101000001010;
10'b0011011110: fsqrtinv_table = 23'b00101110010111110100101;
10'b0011011111: fsqrtinv_table = 23'b00101110001010101001111;
10'b0011100000: fsqrtinv_table = 23'b00101101111101100000110;
10'b0011100001: fsqrtinv_table = 23'b00101101110000011001011;
10'b0011100010: fsqrtinv_table = 23'b00101101100011010011110;
10'b0011100011: fsqrtinv_table = 23'b00101101010110001111110;
10'b0011100100: fsqrtinv_table = 23'b00101101001001001101100;
10'b0011100101: fsqrtinv_table = 23'b00101100111100001100111;
10'b0011100110: fsqrtinv_table = 23'b00101100101111001110000;
10'b0011100111: fsqrtinv_table = 23'b00101100100010010000110;
10'b0011101000: fsqrtinv_table = 23'b00101100010101010101001;
10'b0011101001: fsqrtinv_table = 23'b00101100001000011011010;
10'b0011101010: fsqrtinv_table = 23'b00101011111011100011000;
10'b0011101011: fsqrtinv_table = 23'b00101011101110101100100;
10'b0011101100: fsqrtinv_table = 23'b00101011100001110111100;
10'b0011101101: fsqrtinv_table = 23'b00101011010101000100010;
10'b0011101110: fsqrtinv_table = 23'b00101011001000010010101;
10'b0011101111: fsqrtinv_table = 23'b00101010111011100010101;
10'b0011110000: fsqrtinv_table = 23'b00101010101110110100010;
10'b0011110001: fsqrtinv_table = 23'b00101010100010000111100;
10'b0011110010: fsqrtinv_table = 23'b00101010010101011100011;
10'b0011110011: fsqrtinv_table = 23'b00101010001000110010111;
10'b0011110100: fsqrtinv_table = 23'b00101001111100001010111;
10'b0011110101: fsqrtinv_table = 23'b00101001101111100100101;
10'b0011110110: fsqrtinv_table = 23'b00101001100010111111111;
10'b0011110111: fsqrtinv_table = 23'b00101001010110011100110;
10'b0011111000: fsqrtinv_table = 23'b00101001001001111011001;
10'b0011111001: fsqrtinv_table = 23'b00101000111101011011010;
10'b0011111010: fsqrtinv_table = 23'b00101000110000111100111;
10'b0011111011: fsqrtinv_table = 23'b00101000100100100000000;
10'b0011111100: fsqrtinv_table = 23'b00101000011000000100110;
10'b0011111101: fsqrtinv_table = 23'b00101000001011101011000;
10'b0011111110: fsqrtinv_table = 23'b00100111111111010010111;
10'b0011111111: fsqrtinv_table = 23'b00100111110010111100011;
10'b0100000000: fsqrtinv_table = 23'b00100111100110100111010;
10'b0100000001: fsqrtinv_table = 23'b00100111011010010011110;
10'b0100000010: fsqrtinv_table = 23'b00100111001110000001110;
10'b0100000011: fsqrtinv_table = 23'b00100111000001110001011;
10'b0100000100: fsqrtinv_table = 23'b00100110110101100010011;
10'b0100000101: fsqrtinv_table = 23'b00100110101001010101000;
10'b0100000110: fsqrtinv_table = 23'b00100110011101001001001;
10'b0100000111: fsqrtinv_table = 23'b00100110010000111110110;
10'b0100001000: fsqrtinv_table = 23'b00100110000100110101111;
10'b0100001001: fsqrtinv_table = 23'b00100101111000101110100;
10'b0100001010: fsqrtinv_table = 23'b00100101101100101000101;
10'b0100001011: fsqrtinv_table = 23'b00100101100000100100010;
10'b0100001100: fsqrtinv_table = 23'b00100101010100100001011;
10'b0100001101: fsqrtinv_table = 23'b00100101001000100000000;
10'b0100001110: fsqrtinv_table = 23'b00100100111100100000000;
10'b0100001111: fsqrtinv_table = 23'b00100100110000100001101;
10'b0100010000: fsqrtinv_table = 23'b00100100100100100100101;
10'b0100010001: fsqrtinv_table = 23'b00100100011000101001000;
10'b0100010010: fsqrtinv_table = 23'b00100100001100101111000;
10'b0100010011: fsqrtinv_table = 23'b00100100000000110110011;
10'b0100010100: fsqrtinv_table = 23'b00100011110100111111001;
10'b0100010101: fsqrtinv_table = 23'b00100011101001001001011;
10'b0100010110: fsqrtinv_table = 23'b00100011011101010101001;
10'b0100010111: fsqrtinv_table = 23'b00100011010001100010010;
10'b0100011000: fsqrtinv_table = 23'b00100011000101110000111;
10'b0100011001: fsqrtinv_table = 23'b00100010111010000000111;
10'b0100011010: fsqrtinv_table = 23'b00100010101110010010010;
10'b0100011011: fsqrtinv_table = 23'b00100010100010100101001;
10'b0100011100: fsqrtinv_table = 23'b00100010010110111001010;
10'b0100011101: fsqrtinv_table = 23'b00100010001011001111000;
10'b0100011110: fsqrtinv_table = 23'b00100001111111100110000;
10'b0100011111: fsqrtinv_table = 23'b00100001110011111110100;
10'b0100100000: fsqrtinv_table = 23'b00100001101000011000011;
10'b0100100001: fsqrtinv_table = 23'b00100001011100110011100;
10'b0100100010: fsqrtinv_table = 23'b00100001010001010000001;
10'b0100100011: fsqrtinv_table = 23'b00100001000101101110010;
10'b0100100100: fsqrtinv_table = 23'b00100000111010001101101;
10'b0100100101: fsqrtinv_table = 23'b00100000101110101110011;
10'b0100100110: fsqrtinv_table = 23'b00100000100011010000100;
10'b0100100111: fsqrtinv_table = 23'b00100000010111110100000;
10'b0100101000: fsqrtinv_table = 23'b00100000001100011000110;
10'b0100101001: fsqrtinv_table = 23'b00100000000000111111000;
10'b0100101010: fsqrtinv_table = 23'b00011111110101100110101;
10'b0100101011: fsqrtinv_table = 23'b00011111101010001111100;
10'b0100101100: fsqrtinv_table = 23'b00011111011110111001110;
10'b0100101101: fsqrtinv_table = 23'b00011111010011100101010;
10'b0100101110: fsqrtinv_table = 23'b00011111001000010010010;
10'b0100101111: fsqrtinv_table = 23'b00011110111101000000100;
10'b0100110000: fsqrtinv_table = 23'b00011110110001110000001;
10'b0100110001: fsqrtinv_table = 23'b00011110100110100001000;
10'b0100110010: fsqrtinv_table = 23'b00011110011011010011010;
10'b0100110011: fsqrtinv_table = 23'b00011110010000000110110;
10'b0100110100: fsqrtinv_table = 23'b00011110000100111011101;
10'b0100110101: fsqrtinv_table = 23'b00011101111001110001110;
10'b0100110110: fsqrtinv_table = 23'b00011101101110101001010;
10'b0100110111: fsqrtinv_table = 23'b00011101100011100010000;
10'b0100111000: fsqrtinv_table = 23'b00011101011000011100000;
10'b0100111001: fsqrtinv_table = 23'b00011101001101010111011;
10'b0100111010: fsqrtinv_table = 23'b00011101000010010100000;
10'b0100111011: fsqrtinv_table = 23'b00011100110111010001111;
10'b0100111100: fsqrtinv_table = 23'b00011100101100010001001;
10'b0100111101: fsqrtinv_table = 23'b00011100100001010001101;
10'b0100111110: fsqrtinv_table = 23'b00011100010110010011011;
10'b0100111111: fsqrtinv_table = 23'b00011100001011010110011;
10'b0101000000: fsqrtinv_table = 23'b00011100000000011010101;
10'b0101000001: fsqrtinv_table = 23'b00011011110101100000001;
10'b0101000010: fsqrtinv_table = 23'b00011011101010100111000;
10'b0101000011: fsqrtinv_table = 23'b00011011011111101111000;
10'b0101000100: fsqrtinv_table = 23'b00011011010100111000010;
10'b0101000101: fsqrtinv_table = 23'b00011011001010000010111;
10'b0101000110: fsqrtinv_table = 23'b00011010111111001110101;
10'b0101000111: fsqrtinv_table = 23'b00011010110100011011101;
10'b0101001000: fsqrtinv_table = 23'b00011010101001101001111;
10'b0101001001: fsqrtinv_table = 23'b00011010011110111001011;
10'b0101001010: fsqrtinv_table = 23'b00011010010100001010001;
10'b0101001011: fsqrtinv_table = 23'b00011010001001011100000;
10'b0101001100: fsqrtinv_table = 23'b00011001111110101111001;
10'b0101001101: fsqrtinv_table = 23'b00011001110100000011100;
10'b0101001110: fsqrtinv_table = 23'b00011001101001011001001;
10'b0101001111: fsqrtinv_table = 23'b00011001011110101111111;
10'b0101010000: fsqrtinv_table = 23'b00011001010100000111111;
10'b0101010001: fsqrtinv_table = 23'b00011001001001100001001;
10'b0101010010: fsqrtinv_table = 23'b00011000111110111011100;
10'b0101010011: fsqrtinv_table = 23'b00011000110100010111001;
10'b0101010100: fsqrtinv_table = 23'b00011000101001110011111;
10'b0101010101: fsqrtinv_table = 23'b00011000011111010001111;
10'b0101010110: fsqrtinv_table = 23'b00011000010100110001000;
10'b0101010111: fsqrtinv_table = 23'b00011000001010010001011;
10'b0101011000: fsqrtinv_table = 23'b00010111111111110010111;
10'b0101011001: fsqrtinv_table = 23'b00010111110101010101101;
10'b0101011010: fsqrtinv_table = 23'b00010111101010111001011;
10'b0101011011: fsqrtinv_table = 23'b00010111100000011110100;
10'b0101011100: fsqrtinv_table = 23'b00010111010110000100101;
10'b0101011101: fsqrtinv_table = 23'b00010111001011101100000;
10'b0101011110: fsqrtinv_table = 23'b00010111000001010100100;
10'b0101011111: fsqrtinv_table = 23'b00010110110110111110001;
10'b0101100000: fsqrtinv_table = 23'b00010110101100101001000;
10'b0101100001: fsqrtinv_table = 23'b00010110100010010100111;
10'b0101100010: fsqrtinv_table = 23'b00010110011000000010000;
10'b0101100011: fsqrtinv_table = 23'b00010110001101110000010;
10'b0101100100: fsqrtinv_table = 23'b00010110000011011111101;
10'b0101100101: fsqrtinv_table = 23'b00010101111001010000001;
10'b0101100110: fsqrtinv_table = 23'b00010101101111000001110;
10'b0101100111: fsqrtinv_table = 23'b00010101100100110100100;
10'b0101101000: fsqrtinv_table = 23'b00010101011010101000100;
10'b0101101001: fsqrtinv_table = 23'b00010101010000011101100;
10'b0101101010: fsqrtinv_table = 23'b00010101000110010011101;
10'b0101101011: fsqrtinv_table = 23'b00010100111100001010111;
10'b0101101100: fsqrtinv_table = 23'b00010100110010000011010;
10'b0101101101: fsqrtinv_table = 23'b00010100100111111100101;
10'b0101101110: fsqrtinv_table = 23'b00010100011101110111010;
10'b0101101111: fsqrtinv_table = 23'b00010100010011110010111;
10'b0101110000: fsqrtinv_table = 23'b00010100001001101111101;
10'b0101110001: fsqrtinv_table = 23'b00010011111111101101100;
10'b0101110010: fsqrtinv_table = 23'b00010011110101101100100;
10'b0101110011: fsqrtinv_table = 23'b00010011101011101100100;
10'b0101110100: fsqrtinv_table = 23'b00010011100001101101101;
10'b0101110101: fsqrtinv_table = 23'b00010011010111101111111;
10'b0101110110: fsqrtinv_table = 23'b00010011001101110011010;
10'b0101110111: fsqrtinv_table = 23'b00010011000011110111101;
10'b0101111000: fsqrtinv_table = 23'b00010010111001111101000;
10'b0101111001: fsqrtinv_table = 23'b00010010110000000011100;
10'b0101111010: fsqrtinv_table = 23'b00010010100110001011001;
10'b0101111011: fsqrtinv_table = 23'b00010010011100010011110;
10'b0101111100: fsqrtinv_table = 23'b00010010010010011101100;
10'b0101111101: fsqrtinv_table = 23'b00010010001000101000010;
10'b0101111110: fsqrtinv_table = 23'b00010001111110110100001;
10'b0101111111: fsqrtinv_table = 23'b00010001110101000001000;
10'b0110000000: fsqrtinv_table = 23'b00010001101011001110111;
10'b0110000001: fsqrtinv_table = 23'b00010001100001011101111;
10'b0110000010: fsqrtinv_table = 23'b00010001010111101101111;
10'b0110000011: fsqrtinv_table = 23'b00010001001101111111000;
10'b0110000100: fsqrtinv_table = 23'b00010001000100010001001;
10'b0110000101: fsqrtinv_table = 23'b00010000111010100100010;
10'b0110000110: fsqrtinv_table = 23'b00010000110000111000011;
10'b0110000111: fsqrtinv_table = 23'b00010000100111001101101;
10'b0110001000: fsqrtinv_table = 23'b00010000011101100011110;
10'b0110001001: fsqrtinv_table = 23'b00010000010011111011000;
10'b0110001010: fsqrtinv_table = 23'b00010000001010010011011;
10'b0110001011: fsqrtinv_table = 23'b00010000000000101100101;
10'b0110001100: fsqrtinv_table = 23'b00001111110111000110111;
10'b0110001101: fsqrtinv_table = 23'b00001111101101100010010;
10'b0110001110: fsqrtinv_table = 23'b00001111100011111110101;
10'b0110001111: fsqrtinv_table = 23'b00001111011010011011111;
10'b0110010000: fsqrtinv_table = 23'b00001111010000111010010;
10'b0110010001: fsqrtinv_table = 23'b00001111000111011001101;
10'b0110010010: fsqrtinv_table = 23'b00001110111101111010000;
10'b0110010011: fsqrtinv_table = 23'b00001110110100011011010;
10'b0110010100: fsqrtinv_table = 23'b00001110101010111101101;
10'b0110010101: fsqrtinv_table = 23'b00001110100001100001000;
10'b0110010110: fsqrtinv_table = 23'b00001110011000000101010;
10'b0110010111: fsqrtinv_table = 23'b00001110001110101010101;
10'b0110011000: fsqrtinv_table = 23'b00001110000101010000111;
10'b0110011001: fsqrtinv_table = 23'b00001101111011111000001;
10'b0110011010: fsqrtinv_table = 23'b00001101110010100000011;
10'b0110011011: fsqrtinv_table = 23'b00001101101001001001101;
10'b0110011100: fsqrtinv_table = 23'b00001101011111110011110;
10'b0110011101: fsqrtinv_table = 23'b00001101010110011110111;
10'b0110011110: fsqrtinv_table = 23'b00001101001101001011000;
10'b0110011111: fsqrtinv_table = 23'b00001101000011111000001;
10'b0110100000: fsqrtinv_table = 23'b00001100111010100110010;
10'b0110100001: fsqrtinv_table = 23'b00001100110001010101010;
10'b0110100010: fsqrtinv_table = 23'b00001100101000000101001;
10'b0110100011: fsqrtinv_table = 23'b00001100011110110110001;
10'b0110100100: fsqrtinv_table = 23'b00001100010101101000000;
10'b0110100101: fsqrtinv_table = 23'b00001100001100011010110;
10'b0110100110: fsqrtinv_table = 23'b00001100000011001110100;
10'b0110100111: fsqrtinv_table = 23'b00001011111010000011010;
10'b0110101000: fsqrtinv_table = 23'b00001011110000111000111;
10'b0110101001: fsqrtinv_table = 23'b00001011100111101111100;
10'b0110101010: fsqrtinv_table = 23'b00001011011110100111000;
10'b0110101011: fsqrtinv_table = 23'b00001011010101011111100;
10'b0110101100: fsqrtinv_table = 23'b00001011001100011000111;
10'b0110101101: fsqrtinv_table = 23'b00001011000011010011010;
10'b0110101110: fsqrtinv_table = 23'b00001010111010001110100;
10'b0110101111: fsqrtinv_table = 23'b00001010110001001010101;
10'b0110110000: fsqrtinv_table = 23'b00001010101000000111110;
10'b0110110001: fsqrtinv_table = 23'b00001010011111000101110;
10'b0110110010: fsqrtinv_table = 23'b00001010010110000100101;
10'b0110110011: fsqrtinv_table = 23'b00001010001101000100100;
10'b0110110100: fsqrtinv_table = 23'b00001010000100000101010;
10'b0110110101: fsqrtinv_table = 23'b00001001111011000111000;
10'b0110110110: fsqrtinv_table = 23'b00001001110010001001100;
10'b0110110111: fsqrtinv_table = 23'b00001001101001001101000;
10'b0110111000: fsqrtinv_table = 23'b00001001100000010001011;
10'b0110111001: fsqrtinv_table = 23'b00001001010111010110101;
10'b0110111010: fsqrtinv_table = 23'b00001001001110011100111;
10'b0110111011: fsqrtinv_table = 23'b00001001000101100011111;
10'b0110111100: fsqrtinv_table = 23'b00001000111100101011111;
10'b0110111101: fsqrtinv_table = 23'b00001000110011110100110;
10'b0110111110: fsqrtinv_table = 23'b00001000101010111110100;
10'b0110111111: fsqrtinv_table = 23'b00001000100010001001001;
10'b0111000000: fsqrtinv_table = 23'b00001000011001010100101;
10'b0111000001: fsqrtinv_table = 23'b00001000010000100001000;
10'b0111000010: fsqrtinv_table = 23'b00001000000111101110010;
10'b0111000011: fsqrtinv_table = 23'b00000111111110111100100;
10'b0111000100: fsqrtinv_table = 23'b00000111110110001011100;
10'b0111000101: fsqrtinv_table = 23'b00000111101101011011011;
10'b0111000110: fsqrtinv_table = 23'b00000111100100101100001;
10'b0111000111: fsqrtinv_table = 23'b00000111011011111101110;
10'b0111001000: fsqrtinv_table = 23'b00000111010011010000010;
10'b0111001001: fsqrtinv_table = 23'b00000111001010100011101;
10'b0111001010: fsqrtinv_table = 23'b00000111000001110111111;
10'b0111001011: fsqrtinv_table = 23'b00000110111001001101000;
10'b0111001100: fsqrtinv_table = 23'b00000110110000100010111;
10'b0111001101: fsqrtinv_table = 23'b00000110100111111001110;
10'b0111001110: fsqrtinv_table = 23'b00000110011111010001011;
10'b0111001111: fsqrtinv_table = 23'b00000110010110101001111;
10'b0111010000: fsqrtinv_table = 23'b00000110001110000011010;
10'b0111010001: fsqrtinv_table = 23'b00000110000101011101011;
10'b0111010010: fsqrtinv_table = 23'b00000101111100111000011;
10'b0111010011: fsqrtinv_table = 23'b00000101110100010100010;
10'b0111010100: fsqrtinv_table = 23'b00000101101011110001000;
10'b0111010101: fsqrtinv_table = 23'b00000101100011001110101;
10'b0111010110: fsqrtinv_table = 23'b00000101011010101101000;
10'b0111010111: fsqrtinv_table = 23'b00000101010010001100001;
10'b0111011000: fsqrtinv_table = 23'b00000101001001101100010;
10'b0111011001: fsqrtinv_table = 23'b00000101000001001101001;
10'b0111011010: fsqrtinv_table = 23'b00000100111000101110110;
10'b0111011011: fsqrtinv_table = 23'b00000100110000010001011;
10'b0111011100: fsqrtinv_table = 23'b00000100100111110100110;
10'b0111011101: fsqrtinv_table = 23'b00000100011111011000111;
10'b0111011110: fsqrtinv_table = 23'b00000100010110111101111;
10'b0111011111: fsqrtinv_table = 23'b00000100001110100011101;
10'b0111100000: fsqrtinv_table = 23'b00000100000110001010010;
10'b0111100001: fsqrtinv_table = 23'b00000011111101110001110;
10'b0111100010: fsqrtinv_table = 23'b00000011110101011010000;
10'b0111100011: fsqrtinv_table = 23'b00000011101101000011000;
10'b0111100100: fsqrtinv_table = 23'b00000011100100101100111;
10'b0111100101: fsqrtinv_table = 23'b00000011011100010111100;
10'b0111100110: fsqrtinv_table = 23'b00000011010100000011000;
10'b0111100111: fsqrtinv_table = 23'b00000011001011101111010;
10'b0111101000: fsqrtinv_table = 23'b00000011000011011100010;
10'b0111101001: fsqrtinv_table = 23'b00000010111011001010001;
10'b0111101010: fsqrtinv_table = 23'b00000010110010111000110;
10'b0111101011: fsqrtinv_table = 23'b00000010101010101000010;
10'b0111101100: fsqrtinv_table = 23'b00000010100010011000100;
10'b0111101101: fsqrtinv_table = 23'b00000010011010001001100;
10'b0111101110: fsqrtinv_table = 23'b00000010010001111011010;
10'b0111101111: fsqrtinv_table = 23'b00000010001001101101111;
10'b0111110000: fsqrtinv_table = 23'b00000010000001100001010;
10'b0111110001: fsqrtinv_table = 23'b00000001111001010101011;
10'b0111110010: fsqrtinv_table = 23'b00000001110001001010011;
10'b0111110011: fsqrtinv_table = 23'b00000001101001000000000;
10'b0111110100: fsqrtinv_table = 23'b00000001100000110110100;
10'b0111110101: fsqrtinv_table = 23'b00000001011000101101110;
10'b0111110110: fsqrtinv_table = 23'b00000001010000100101110;
10'b0111110111: fsqrtinv_table = 23'b00000001001000011110101;
10'b0111111000: fsqrtinv_table = 23'b00000001000000011000001;
10'b0111111001: fsqrtinv_table = 23'b00000000111000010010100;
10'b0111111010: fsqrtinv_table = 23'b00000000110000001101101;
10'b0111111011: fsqrtinv_table = 23'b00000000101000001001011;
10'b0111111100: fsqrtinv_table = 23'b00000000100000000110000;
10'b0111111101: fsqrtinv_table = 23'b00000000011000000011011;
10'b0111111110: fsqrtinv_table = 23'b00000000010000000001100;
10'b0111111111: fsqrtinv_table = 23'b00000000001000000000011;
10'b1000000000: fsqrtinv_table = 23'b00000000000000000000000;
10'b1000000001: fsqrtinv_table = 23'b11111111100000000011000;
10'b1000000010: fsqrtinv_table = 23'b11111111000000001100000;
10'b1000000011: fsqrtinv_table = 23'b11111110100000011010111;
10'b1000000100: fsqrtinv_table = 23'b11111110000000101111110;
10'b1000000101: fsqrtinv_table = 23'b11111101100001001010011;
10'b1000000110: fsqrtinv_table = 23'b11111101000001101011000;
10'b1000000111: fsqrtinv_table = 23'b11111100100010010001011;
10'b1000001000: fsqrtinv_table = 23'b11111100000010111101100;
10'b1000001001: fsqrtinv_table = 23'b11111011100011101111100;
10'b1000001010: fsqrtinv_table = 23'b11111011000100100111010;
10'b1000001011: fsqrtinv_table = 23'b11111010100101100100101;
10'b1000001100: fsqrtinv_table = 23'b11111010000110100111110;
10'b1000001101: fsqrtinv_table = 23'b11111001100111110000100;
10'b1000001110: fsqrtinv_table = 23'b11111001001000111110111;
10'b1000001111: fsqrtinv_table = 23'b11111000101010010010111;
10'b1000010000: fsqrtinv_table = 23'b11111000001011101100100;
10'b1000010001: fsqrtinv_table = 23'b11110111101101001011101;
10'b1000010010: fsqrtinv_table = 23'b11110111001110110000011;
10'b1000010011: fsqrtinv_table = 23'b11110110110000011010100;
10'b1000010100: fsqrtinv_table = 23'b11110110010010001010010;
10'b1000010101: fsqrtinv_table = 23'b11110101110011111111011;
10'b1000010110: fsqrtinv_table = 23'b11110101010101111001111;
10'b1000010111: fsqrtinv_table = 23'b11110100110111111001111;
10'b1000011000: fsqrtinv_table = 23'b11110100011001111111001;
10'b1000011001: fsqrtinv_table = 23'b11110011111100001001111;
10'b1000011010: fsqrtinv_table = 23'b11110011011110011001111;
10'b1000011011: fsqrtinv_table = 23'b11110011000000101111001;
10'b1000011100: fsqrtinv_table = 23'b11110010100011001001110;
10'b1000011101: fsqrtinv_table = 23'b11110010000101101001100;
10'b1000011110: fsqrtinv_table = 23'b11110001101000001110101;
10'b1000011111: fsqrtinv_table = 23'b11110001001010111000111;
10'b1000100000: fsqrtinv_table = 23'b11110000101101101000010;
10'b1000100001: fsqrtinv_table = 23'b11110000010000011100111;
10'b1000100010: fsqrtinv_table = 23'b11101111110011010110101;
10'b1000100011: fsqrtinv_table = 23'b11101111010110010101100;
10'b1000100100: fsqrtinv_table = 23'b11101110111001011001011;
10'b1000100101: fsqrtinv_table = 23'b11101110011100100010011;
10'b1000100110: fsqrtinv_table = 23'b11101101111111110000011;
10'b1000100111: fsqrtinv_table = 23'b11101101100011000011011;
10'b1000101000: fsqrtinv_table = 23'b11101101000110011011100;
10'b1000101001: fsqrtinv_table = 23'b11101100101001111000100;
10'b1000101010: fsqrtinv_table = 23'b11101100001101011010011;
10'b1000101011: fsqrtinv_table = 23'b11101011110001000001010;
10'b1000101100: fsqrtinv_table = 23'b11101011010100101101001;
10'b1000101101: fsqrtinv_table = 23'b11101010111000011101110;
10'b1000101110: fsqrtinv_table = 23'b11101010011100010011010;
10'b1000101111: fsqrtinv_table = 23'b11101010000000001101101;
10'b1000110000: fsqrtinv_table = 23'b11101001100100001100111;
10'b1000110001: fsqrtinv_table = 23'b11101001001000010000111;
10'b1000110010: fsqrtinv_table = 23'b11101000101100011001101;
10'b1000110011: fsqrtinv_table = 23'b11101000010000100111001;
10'b1000110100: fsqrtinv_table = 23'b11100111110100111001011;
10'b1000110101: fsqrtinv_table = 23'b11100111011001010000010;
10'b1000110110: fsqrtinv_table = 23'b11100110111101101100000;
10'b1000110111: fsqrtinv_table = 23'b11100110100010001100010;
10'b1000111000: fsqrtinv_table = 23'b11100110000110110001010;
10'b1000111001: fsqrtinv_table = 23'b11100101101011011010111;
10'b1000111010: fsqrtinv_table = 23'b11100101010000001001000;
10'b1000111011: fsqrtinv_table = 23'b11100100110100111011110;
10'b1000111100: fsqrtinv_table = 23'b11100100011001110011001;
10'b1000111101: fsqrtinv_table = 23'b11100011111110101111001;
10'b1000111110: fsqrtinv_table = 23'b11100011100011101111100;
10'b1000111111: fsqrtinv_table = 23'b11100011001000110100011;
10'b1001000000: fsqrtinv_table = 23'b11100010101101111101111;
10'b1001000001: fsqrtinv_table = 23'b11100010010011001011110;
10'b1001000010: fsqrtinv_table = 23'b11100001111000011110001;
10'b1001000011: fsqrtinv_table = 23'b11100001011101110100111;
10'b1001000100: fsqrtinv_table = 23'b11100001000011010000001;
10'b1001000101: fsqrtinv_table = 23'b11100000101000101111101;
10'b1001000110: fsqrtinv_table = 23'b11100000001110010011101;
10'b1001000111: fsqrtinv_table = 23'b11011111110011111100000;
10'b1001001000: fsqrtinv_table = 23'b11011111011001101000101;
10'b1001001001: fsqrtinv_table = 23'b11011110111111011001101;
10'b1001001010: fsqrtinv_table = 23'b11011110100101001110111;
10'b1001001011: fsqrtinv_table = 23'b11011110001011001000011;
10'b1001001100: fsqrtinv_table = 23'b11011101110001000110010;
10'b1001001101: fsqrtinv_table = 23'b11011101010111001000010;
10'b1001001110: fsqrtinv_table = 23'b11011100111101001110100;
10'b1001001111: fsqrtinv_table = 23'b11011100100011011001000;
10'b1001010000: fsqrtinv_table = 23'b11011100001001100111110;
10'b1001010001: fsqrtinv_table = 23'b11011011101111111010101;
10'b1001010010: fsqrtinv_table = 23'b11011011010110010001101;
10'b1001010011: fsqrtinv_table = 23'b11011010111100101100110;
10'b1001010100: fsqrtinv_table = 23'b11011010100011001100000;
10'b1001010101: fsqrtinv_table = 23'b11011010001001101111100;
10'b1001010110: fsqrtinv_table = 23'b11011001110000010110111;
10'b1001010111: fsqrtinv_table = 23'b11011001010111000010100;
10'b1001011000: fsqrtinv_table = 23'b11011000111101110010000;
10'b1001011001: fsqrtinv_table = 23'b11011000100100100101101;
10'b1001011010: fsqrtinv_table = 23'b11011000001011011101010;
10'b1001011011: fsqrtinv_table = 23'b11010111110010011001000;
10'b1001011100: fsqrtinv_table = 23'b11010111011001011000101;
10'b1001011101: fsqrtinv_table = 23'b11010111000000011100010;
10'b1001011110: fsqrtinv_table = 23'b11010110100111100011110;
10'b1001011111: fsqrtinv_table = 23'b11010110001110101111010;
10'b1001100000: fsqrtinv_table = 23'b11010101110101111110101;
10'b1001100001: fsqrtinv_table = 23'b11010101011101010010000;
10'b1001100010: fsqrtinv_table = 23'b11010101000100101001001;
10'b1001100011: fsqrtinv_table = 23'b11010100101100000100010;
10'b1001100100: fsqrtinv_table = 23'b11010100010011100011010;
10'b1001100101: fsqrtinv_table = 23'b11010011111011000110000;
10'b1001100110: fsqrtinv_table = 23'b11010011100010101100101;
10'b1001100111: fsqrtinv_table = 23'b11010011001010010111000;
10'b1001101000: fsqrtinv_table = 23'b11010010110010000101010;
10'b1001101001: fsqrtinv_table = 23'b11010010011001110111010;
10'b1001101010: fsqrtinv_table = 23'b11010010000001101101000;
10'b1001101011: fsqrtinv_table = 23'b11010001101001100110100;
10'b1001101100: fsqrtinv_table = 23'b11010001010001100011101;
10'b1001101101: fsqrtinv_table = 23'b11010000111001100100101;
10'b1001101110: fsqrtinv_table = 23'b11010000100001101001010;
10'b1001101111: fsqrtinv_table = 23'b11010000001001110001101;
10'b1001110000: fsqrtinv_table = 23'b11001111110001111101101;
10'b1001110001: fsqrtinv_table = 23'b11001111011010001101010;
10'b1001110010: fsqrtinv_table = 23'b11001111000010100000101;
10'b1001110011: fsqrtinv_table = 23'b11001110101010110111101;
10'b1001110100: fsqrtinv_table = 23'b11001110010011010010001;
10'b1001110101: fsqrtinv_table = 23'b11001101111011110000010;
10'b1001110110: fsqrtinv_table = 23'b11001101100100010010001;
10'b1001110111: fsqrtinv_table = 23'b11001101001100110111011;
10'b1001111000: fsqrtinv_table = 23'b11001100110101100000010;
10'b1001111001: fsqrtinv_table = 23'b11001100011110001100110;
10'b1001111010: fsqrtinv_table = 23'b11001100000110111100101;
10'b1001111011: fsqrtinv_table = 23'b11001011101111110000001;
10'b1001111100: fsqrtinv_table = 23'b11001011011000100111001;
10'b1001111101: fsqrtinv_table = 23'b11001011000001100001101;
10'b1001111110: fsqrtinv_table = 23'b11001010101010011111100;
10'b1001111111: fsqrtinv_table = 23'b11001010010011100000111;
10'b1010000000: fsqrtinv_table = 23'b11001001111100100101110;
10'b1010000001: fsqrtinv_table = 23'b11001001100101101110000;
10'b1010000010: fsqrtinv_table = 23'b11001001001110111001110;
10'b1010000011: fsqrtinv_table = 23'b11001000111000001000111;
10'b1010000100: fsqrtinv_table = 23'b11001000100001011011011;
10'b1010000101: fsqrtinv_table = 23'b11001000001010110001010;
10'b1010000110: fsqrtinv_table = 23'b11000111110100001010100;
10'b1010000111: fsqrtinv_table = 23'b11000111011101100111001;
10'b1010001000: fsqrtinv_table = 23'b11000111000111000111001;
10'b1010001001: fsqrtinv_table = 23'b11000110110000101010011;
10'b1010001010: fsqrtinv_table = 23'b11000110011010010001000;
10'b1010001011: fsqrtinv_table = 23'b11000110000011111010111;
10'b1010001100: fsqrtinv_table = 23'b11000101101101101000001;
10'b1010001101: fsqrtinv_table = 23'b11000101010111011000101;
10'b1010001110: fsqrtinv_table = 23'b11000101000001001100011;
10'b1010001111: fsqrtinv_table = 23'b11000100101011000011011;
10'b1010010000: fsqrtinv_table = 23'b11000100010100111101101;
10'b1010010001: fsqrtinv_table = 23'b11000011111110111011000;
10'b1010010010: fsqrtinv_table = 23'b11000011101000111011110;
10'b1010010011: fsqrtinv_table = 23'b11000011010010111111101;
10'b1010010100: fsqrtinv_table = 23'b11000010111101000110110;
10'b1010010101: fsqrtinv_table = 23'b11000010100111010001000;
10'b1010010110: fsqrtinv_table = 23'b11000010010001011110011;
10'b1010010111: fsqrtinv_table = 23'b11000001111011101111000;
10'b1010011000: fsqrtinv_table = 23'b11000001100110000010110;
10'b1010011001: fsqrtinv_table = 23'b11000001010000011001100;
10'b1010011010: fsqrtinv_table = 23'b11000000111010110011100;
10'b1010011011: fsqrtinv_table = 23'b11000000100101010000101;
10'b1010011100: fsqrtinv_table = 23'b11000000001111110000111;
10'b1010011101: fsqrtinv_table = 23'b10111111111010010100001;
10'b1010011110: fsqrtinv_table = 23'b10111111100100111010100;
10'b1010011111: fsqrtinv_table = 23'b10111111001111100011111;
10'b1010100000: fsqrtinv_table = 23'b10111110111010010000011;
10'b1010100001: fsqrtinv_table = 23'b10111110100100111111111;
10'b1010100010: fsqrtinv_table = 23'b10111110001111110010011;
10'b1010100011: fsqrtinv_table = 23'b10111101111010100111111;
10'b1010100100: fsqrtinv_table = 23'b10111101100101100000100;
10'b1010100101: fsqrtinv_table = 23'b10111101010000011100000;
10'b1010100110: fsqrtinv_table = 23'b10111100111011011010101;
10'b1010100111: fsqrtinv_table = 23'b10111100100110011100001;
10'b1010101000: fsqrtinv_table = 23'b10111100010001100000101;
10'b1010101001: fsqrtinv_table = 23'b10111011111100101000000;
10'b1010101010: fsqrtinv_table = 23'b10111011100111110010011;
10'b1010101011: fsqrtinv_table = 23'b10111011010010111111101;
10'b1010101100: fsqrtinv_table = 23'b10111010111110001111111;
10'b1010101101: fsqrtinv_table = 23'b10111010101001100011000;
10'b1010101110: fsqrtinv_table = 23'b10111010010100111001000;
10'b1010101111: fsqrtinv_table = 23'b10111010000000010010000;
10'b1010110000: fsqrtinv_table = 23'b10111001101011101101110;
10'b1010110001: fsqrtinv_table = 23'b10111001010111001100011;
10'b1010110010: fsqrtinv_table = 23'b10111001000010101101111;
10'b1010110011: fsqrtinv_table = 23'b10111000101110010010010;
10'b1010110100: fsqrtinv_table = 23'b10111000011001111001100;
10'b1010110101: fsqrtinv_table = 23'b10111000000101100011100;
10'b1010110110: fsqrtinv_table = 23'b10110111110001010000010;
10'b1010110111: fsqrtinv_table = 23'b10110111011100111111111;
10'b1010111000: fsqrtinv_table = 23'b10110111001000110010011;
10'b1010111001: fsqrtinv_table = 23'b10110110110100100111101;
10'b1010111010: fsqrtinv_table = 23'b10110110100000011111101;
10'b1010111011: fsqrtinv_table = 23'b10110110001100011010011;
10'b1010111100: fsqrtinv_table = 23'b10110101111000010111111;
10'b1010111101: fsqrtinv_table = 23'b10110101100100011000001;
10'b1010111110: fsqrtinv_table = 23'b10110101010000011011001;
10'b1010111111: fsqrtinv_table = 23'b10110100111100100000110;
10'b1011000000: fsqrtinv_table = 23'b10110100101000101001010;
10'b1011000001: fsqrtinv_table = 23'b10110100010100110100011;
10'b1011000010: fsqrtinv_table = 23'b10110100000001000010010;
10'b1011000011: fsqrtinv_table = 23'b10110011101101010010110;
10'b1011000100: fsqrtinv_table = 23'b10110011011001100110000;
10'b1011000101: fsqrtinv_table = 23'b10110011000101111011110;
10'b1011000110: fsqrtinv_table = 23'b10110010110010010100011;
10'b1011000111: fsqrtinv_table = 23'b10110010011110101111100;
10'b1011001000: fsqrtinv_table = 23'b10110010001011001101011;
10'b1011001001: fsqrtinv_table = 23'b10110001110111101101110;
10'b1011001010: fsqrtinv_table = 23'b10110001100100010000111;
10'b1011001011: fsqrtinv_table = 23'b10110001010000110110100;
10'b1011001100: fsqrtinv_table = 23'b10110000111101011110111;
10'b1011001101: fsqrtinv_table = 23'b10110000101010001001110;
10'b1011001110: fsqrtinv_table = 23'b10110000010110110111010;
10'b1011001111: fsqrtinv_table = 23'b10110000000011100111010;
10'b1011010000: fsqrtinv_table = 23'b10101111110000011001111;
10'b1011010001: fsqrtinv_table = 23'b10101111011101001111000;
10'b1011010010: fsqrtinv_table = 23'b10101111001010000110110;
10'b1011010011: fsqrtinv_table = 23'b10101110110111000001000;
10'b1011010100: fsqrtinv_table = 23'b10101110100011111101110;
10'b1011010101: fsqrtinv_table = 23'b10101110010000111101001;
10'b1011010110: fsqrtinv_table = 23'b10101101111101111111000;
10'b1011010111: fsqrtinv_table = 23'b10101101101011000011010;
10'b1011011000: fsqrtinv_table = 23'b10101101011000001010001;
10'b1011011001: fsqrtinv_table = 23'b10101101000101010011011;
10'b1011011010: fsqrtinv_table = 23'b10101100110010011111010;
10'b1011011011: fsqrtinv_table = 23'b10101100011111101101100;
10'b1011011100: fsqrtinv_table = 23'b10101100001100111110010;
10'b1011011101: fsqrtinv_table = 23'b10101011111010010001100;
10'b1011011110: fsqrtinv_table = 23'b10101011100111100111001;
10'b1011011111: fsqrtinv_table = 23'b10101011010100111111001;
10'b1011100000: fsqrtinv_table = 23'b10101011000010011001101;
10'b1011100001: fsqrtinv_table = 23'b10101010101111110110101;
10'b1011100010: fsqrtinv_table = 23'b10101010011101010110000;
10'b1011100011: fsqrtinv_table = 23'b10101010001010110111110;
10'b1011100100: fsqrtinv_table = 23'b10101001111000011011111;
10'b1011100101: fsqrtinv_table = 23'b10101001100110000010011;
10'b1011100110: fsqrtinv_table = 23'b10101001010011101011010;
10'b1011100111: fsqrtinv_table = 23'b10101001000001010110101;
10'b1011101000: fsqrtinv_table = 23'b10101000101111000100010;
10'b1011101001: fsqrtinv_table = 23'b10101000011100110100010;
10'b1011101010: fsqrtinv_table = 23'b10101000001010100110101;
10'b1011101011: fsqrtinv_table = 23'b10100111111000011011011;
10'b1011101100: fsqrtinv_table = 23'b10100111100110010010011;
10'b1011101101: fsqrtinv_table = 23'b10100111010100001011110;
10'b1011101110: fsqrtinv_table = 23'b10100111000010000111011;
10'b1011101111: fsqrtinv_table = 23'b10100110110000000101011;
10'b1011110000: fsqrtinv_table = 23'b10100110011110000101110;
10'b1011110001: fsqrtinv_table = 23'b10100110001100001000010;
10'b1011110010: fsqrtinv_table = 23'b10100101111010001101001;
10'b1011110011: fsqrtinv_table = 23'b10100101101000010100011;
10'b1011110100: fsqrtinv_table = 23'b10100101010110011101110;
10'b1011110101: fsqrtinv_table = 23'b10100101000100101001100;
10'b1011110110: fsqrtinv_table = 23'b10100100110010110111011;
10'b1011110111: fsqrtinv_table = 23'b10100100100001000111101;
10'b1011111000: fsqrtinv_table = 23'b10100100001111011010000;
10'b1011111001: fsqrtinv_table = 23'b10100011111101101110110;
10'b1011111010: fsqrtinv_table = 23'b10100011101100000101101;
10'b1011111011: fsqrtinv_table = 23'b10100011011010011110110;
10'b1011111100: fsqrtinv_table = 23'b10100011001000111010001;
10'b1011111101: fsqrtinv_table = 23'b10100010110111010111101;
10'b1011111110: fsqrtinv_table = 23'b10100010100101110111011;
10'b1011111111: fsqrtinv_table = 23'b10100010010100011001011;
10'b1100000000: fsqrtinv_table = 23'b10100010000010111101100;
10'b1100000001: fsqrtinv_table = 23'b10100001110001100011110;
10'b1100000010: fsqrtinv_table = 23'b10100001100000001100010;
10'b1100000011: fsqrtinv_table = 23'b10100001001110110110111;
10'b1100000100: fsqrtinv_table = 23'b10100000111101100011101;
10'b1100000101: fsqrtinv_table = 23'b10100000101100010010100;
10'b1100000110: fsqrtinv_table = 23'b10100000011011000011101;
10'b1100000111: fsqrtinv_table = 23'b10100000001001110110111;
10'b1100001000: fsqrtinv_table = 23'b10011111111000101100010;
10'b1100001001: fsqrtinv_table = 23'b10011111100111100011101;
10'b1100001010: fsqrtinv_table = 23'b10011111010110011101010;
10'b1100001011: fsqrtinv_table = 23'b10011111000101011000111;
10'b1100001100: fsqrtinv_table = 23'b10011110110100010110110;
10'b1100001101: fsqrtinv_table = 23'b10011110100011010110101;
10'b1100001110: fsqrtinv_table = 23'b10011110010010011000101;
10'b1100001111: fsqrtinv_table = 23'b10011110000001011100101;
10'b1100010000: fsqrtinv_table = 23'b10011101110000100010110;
10'b1100010001: fsqrtinv_table = 23'b10011101011111101011000;
10'b1100010010: fsqrtinv_table = 23'b10011101001110110101010;
10'b1100010011: fsqrtinv_table = 23'b10011100111110000001100;
10'b1100010100: fsqrtinv_table = 23'b10011100101101001111111;
10'b1100010101: fsqrtinv_table = 23'b10011100011100100000010;
10'b1100010110: fsqrtinv_table = 23'b10011100001011110010110;
10'b1100010111: fsqrtinv_table = 23'b10011011111011000111001;
10'b1100011000: fsqrtinv_table = 23'b10011011101010011101101;
10'b1100011001: fsqrtinv_table = 23'b10011011011001110110001;
10'b1100011010: fsqrtinv_table = 23'b10011011001001010000101;
10'b1100011011: fsqrtinv_table = 23'b10011010111000101101001;
10'b1100011100: fsqrtinv_table = 23'b10011010101000001011110;
10'b1100011101: fsqrtinv_table = 23'b10011010010111101100010;
10'b1100011110: fsqrtinv_table = 23'b10011010000111001110110;
10'b1100011111: fsqrtinv_table = 23'b10011001110110110011001;
10'b1100100000: fsqrtinv_table = 23'b10011001100110011001101;
10'b1100100001: fsqrtinv_table = 23'b10011001010110000010000;
10'b1100100010: fsqrtinv_table = 23'b10011001000101101100011;
10'b1100100011: fsqrtinv_table = 23'b10011000110101011000110;
10'b1100100100: fsqrtinv_table = 23'b10011000100101000111000;
10'b1100100101: fsqrtinv_table = 23'b10011000010100110111001;
10'b1100100110: fsqrtinv_table = 23'b10011000000100101001011;
10'b1100100111: fsqrtinv_table = 23'b10010111110100011101011;
10'b1100101000: fsqrtinv_table = 23'b10010111100100010011011;
10'b1100101001: fsqrtinv_table = 23'b10010111010100001011010;
10'b1100101010: fsqrtinv_table = 23'b10010111000100000101001;
10'b1100101011: fsqrtinv_table = 23'b10010110110100000000111;
10'b1100101100: fsqrtinv_table = 23'b10010110100011111110100;
10'b1100101101: fsqrtinv_table = 23'b10010110010011111110000;
10'b1100101110: fsqrtinv_table = 23'b10010110000011111111100;
10'b1100101111: fsqrtinv_table = 23'b10010101110100000010110;
10'b1100110000: fsqrtinv_table = 23'b10010101100100000111111;
10'b1100110001: fsqrtinv_table = 23'b10010101010100001111000;
10'b1100110010: fsqrtinv_table = 23'b10010101000100010111111;
10'b1100110011: fsqrtinv_table = 23'b10010100110100100010101;
10'b1100110100: fsqrtinv_table = 23'b10010100100100101111010;
10'b1100110101: fsqrtinv_table = 23'b10010100010100111101110;
10'b1100110110: fsqrtinv_table = 23'b10010100000101001110001;
10'b1100110111: fsqrtinv_table = 23'b10010011110101100000010;
10'b1100111000: fsqrtinv_table = 23'b10010011100101110100010;
10'b1100111001: fsqrtinv_table = 23'b10010011010110001010000;
10'b1100111010: fsqrtinv_table = 23'b10010011000110100001101;
10'b1100111011: fsqrtinv_table = 23'b10010010110110111011001;
10'b1100111100: fsqrtinv_table = 23'b10010010100111010110011;
10'b1100111101: fsqrtinv_table = 23'b10010010010111110011011;
10'b1100111110: fsqrtinv_table = 23'b10010010001000010010010;
10'b1100111111: fsqrtinv_table = 23'b10010001111000110011000;
10'b1101000000: fsqrtinv_table = 23'b10010001101001010101011;
10'b1101000001: fsqrtinv_table = 23'b10010001011001111001101;
10'b1101000010: fsqrtinv_table = 23'b10010001001010011111101;
10'b1101000011: fsqrtinv_table = 23'b10010000111011000111011;
10'b1101000100: fsqrtinv_table = 23'b10010000101011110000111;
10'b1101000101: fsqrtinv_table = 23'b10010000011100011100010;
10'b1101000110: fsqrtinv_table = 23'b10010000001101001001010;
10'b1101000111: fsqrtinv_table = 23'b10001111111101111000001;
10'b1101001000: fsqrtinv_table = 23'b10001111101110101000101;
10'b1101001001: fsqrtinv_table = 23'b10001111011111011010111;
10'b1101001010: fsqrtinv_table = 23'b10001111010000001111000;
10'b1101001011: fsqrtinv_table = 23'b10001111000001000100110;
10'b1101001100: fsqrtinv_table = 23'b10001110110001111100010;
10'b1101001101: fsqrtinv_table = 23'b10001110100010110101011;
10'b1101001110: fsqrtinv_table = 23'b10001110010011110000011;
10'b1101001111: fsqrtinv_table = 23'b10001110000100101101000;
10'b1101010000: fsqrtinv_table = 23'b10001101110101101011010;
10'b1101010001: fsqrtinv_table = 23'b10001101100110101011010;
10'b1101010010: fsqrtinv_table = 23'b10001101010111101101000;
10'b1101010011: fsqrtinv_table = 23'b10001101001000110000100;
10'b1101010100: fsqrtinv_table = 23'b10001100111001110101100;
10'b1101010101: fsqrtinv_table = 23'b10001100101010111100011;
10'b1101010110: fsqrtinv_table = 23'b10001100011100000100110;
10'b1101010111: fsqrtinv_table = 23'b10001100001101001110111;
10'b1101011000: fsqrtinv_table = 23'b10001011111110011010110;
10'b1101011001: fsqrtinv_table = 23'b10001011101111101000001;
10'b1101011010: fsqrtinv_table = 23'b10001011100000110111010;
10'b1101011011: fsqrtinv_table = 23'b10001011010010001000000;
10'b1101011100: fsqrtinv_table = 23'b10001011000011011010011;
10'b1101011101: fsqrtinv_table = 23'b10001010110100101110100;
10'b1101011110: fsqrtinv_table = 23'b10001010100110000100001;
10'b1101011111: fsqrtinv_table = 23'b10001010010111011011011;
10'b1101100000: fsqrtinv_table = 23'b10001010001000110100011;
10'b1101100001: fsqrtinv_table = 23'b10001001111010001110111;
10'b1101100010: fsqrtinv_table = 23'b10001001101011101011001;
10'b1101100011: fsqrtinv_table = 23'b10001001011101001000111;
10'b1101100100: fsqrtinv_table = 23'b10001001001110101000010;
10'b1101100101: fsqrtinv_table = 23'b10001001000000001001010;
10'b1101100110: fsqrtinv_table = 23'b10001000110001101011111;
10'b1101100111: fsqrtinv_table = 23'b10001000100011010000001;
10'b1101101000: fsqrtinv_table = 23'b10001000010100110101111;
10'b1101101001: fsqrtinv_table = 23'b10001000000110011101010;
10'b1101101010: fsqrtinv_table = 23'b10000111111000000110001;
10'b1101101011: fsqrtinv_table = 23'b10000111101001110000101;
10'b1101101100: fsqrtinv_table = 23'b10000111011011011100110;
10'b1101101101: fsqrtinv_table = 23'b10000111001101001010100;
10'b1101101110: fsqrtinv_table = 23'b10000110111110111001101;
10'b1101101111: fsqrtinv_table = 23'b10000110110000101010100;
10'b1101110000: fsqrtinv_table = 23'b10000110100010011100110;
10'b1101110001: fsqrtinv_table = 23'b10000110010100010000101;
10'b1101110010: fsqrtinv_table = 23'b10000110000110000110001;
10'b1101110011: fsqrtinv_table = 23'b10000101110111111101001;
10'b1101110100: fsqrtinv_table = 23'b10000101101001110101101;
10'b1101110101: fsqrtinv_table = 23'b10000101011011101111101;
10'b1101110110: fsqrtinv_table = 23'b10000101001101101011001;
10'b1101110111: fsqrtinv_table = 23'b10000100111111101000010;
10'b1101111000: fsqrtinv_table = 23'b10000100110001100110111;
10'b1101111001: fsqrtinv_table = 23'b10000100100011100111000;
10'b1101111010: fsqrtinv_table = 23'b10000100010101101000101;
10'b1101111011: fsqrtinv_table = 23'b10000100000111101011110;
10'b1101111100: fsqrtinv_table = 23'b10000011111001110000011;
10'b1101111101: fsqrtinv_table = 23'b10000011101011110110100;
10'b1101111110: fsqrtinv_table = 23'b10000011011101111110001;
10'b1101111111: fsqrtinv_table = 23'b10000011010000000111010;
10'b1110000000: fsqrtinv_table = 23'b10000011000010010001111;
10'b1110000001: fsqrtinv_table = 23'b10000010110100011110000;
10'b1110000010: fsqrtinv_table = 23'b10000010100110101011100;
10'b1110000011: fsqrtinv_table = 23'b10000010011000111010101;
10'b1110000100: fsqrtinv_table = 23'b10000010001011001011001;
10'b1110000101: fsqrtinv_table = 23'b10000001111101011101001;
10'b1110000110: fsqrtinv_table = 23'b10000001101111110000100;
10'b1110000111: fsqrtinv_table = 23'b10000001100010000101011;
10'b1110001000: fsqrtinv_table = 23'b10000001010100011011110;
10'b1110001001: fsqrtinv_table = 23'b10000001000110110011100;
10'b1110001010: fsqrtinv_table = 23'b10000000111001001100110;
10'b1110001011: fsqrtinv_table = 23'b10000000101011100111011;
10'b1110001100: fsqrtinv_table = 23'b10000000011110000011100;
10'b1110001101: fsqrtinv_table = 23'b10000000010000100001001;
10'b1110001110: fsqrtinv_table = 23'b10000000000011000000000;
10'b1110001111: fsqrtinv_table = 23'b01111111110101100000011;
10'b1110010000: fsqrtinv_table = 23'b01111111101000000010010;
10'b1110010001: fsqrtinv_table = 23'b01111111011010100101100;
10'b1110010010: fsqrtinv_table = 23'b01111111001101001010001;
10'b1110010011: fsqrtinv_table = 23'b01111110111111110000001;
10'b1110010100: fsqrtinv_table = 23'b01111110110010010111101;
10'b1110010101: fsqrtinv_table = 23'b01111110100101000000100;
10'b1110010110: fsqrtinv_table = 23'b01111110010111101010110;
10'b1110010111: fsqrtinv_table = 23'b01111110001010010110011;
10'b1110011000: fsqrtinv_table = 23'b01111101111101000011100;
10'b1110011001: fsqrtinv_table = 23'b01111101101111110001111;
10'b1110011010: fsqrtinv_table = 23'b01111101100010100001110;
10'b1110011011: fsqrtinv_table = 23'b01111101010101010010111;
10'b1110011100: fsqrtinv_table = 23'b01111101001000000101100;
10'b1110011101: fsqrtinv_table = 23'b01111100111010111001011;
10'b1110011110: fsqrtinv_table = 23'b01111100101101101110110;
10'b1110011111: fsqrtinv_table = 23'b01111100100000100101011;
10'b1110100000: fsqrtinv_table = 23'b01111100010011011101011;
10'b1110100001: fsqrtinv_table = 23'b01111100000110010110110;
10'b1110100010: fsqrtinv_table = 23'b01111011111001010001100;
10'b1110100011: fsqrtinv_table = 23'b01111011101100001101101;
10'b1110100100: fsqrtinv_table = 23'b01111011011111001011000;
10'b1110100101: fsqrtinv_table = 23'b01111011010010001001111;
10'b1110100110: fsqrtinv_table = 23'b01111011000101001001111;
10'b1110100111: fsqrtinv_table = 23'b01111010111000001011011;
10'b1110101000: fsqrtinv_table = 23'b01111010101011001110001;
10'b1110101001: fsqrtinv_table = 23'b01111010011110010010010;
10'b1110101010: fsqrtinv_table = 23'b01111010010001010111110;
10'b1110101011: fsqrtinv_table = 23'b01111010000100011110100;
10'b1110101100: fsqrtinv_table = 23'b01111001110111100110100;
10'b1110101101: fsqrtinv_table = 23'b01111001101010101111111;
10'b1110101110: fsqrtinv_table = 23'b01111001011101111010101;
10'b1110101111: fsqrtinv_table = 23'b01111001010001000110101;
10'b1110110000: fsqrtinv_table = 23'b01111001000100010011111;
10'b1110110001: fsqrtinv_table = 23'b01111000110111100010100;
10'b1110110010: fsqrtinv_table = 23'b01111000101010110010011;
10'b1110110011: fsqrtinv_table = 23'b01111000011110000011101;
10'b1110110100: fsqrtinv_table = 23'b01111000010001010110001;
10'b1110110101: fsqrtinv_table = 23'b01111000000100101001111;
10'b1110110110: fsqrtinv_table = 23'b01110111110111111110111;
10'b1110110111: fsqrtinv_table = 23'b01110111101011010101010;
10'b1110111000: fsqrtinv_table = 23'b01110111011110101100111;
10'b1110111001: fsqrtinv_table = 23'b01110111010010000101110;
10'b1110111010: fsqrtinv_table = 23'b01110111000101011111111;
10'b1110111011: fsqrtinv_table = 23'b01110110111000111011011;
10'b1110111100: fsqrtinv_table = 23'b01110110101100011000000;
10'b1110111101: fsqrtinv_table = 23'b01110110011111110101111;
10'b1110111110: fsqrtinv_table = 23'b01110110010011010101001;
10'b1110111111: fsqrtinv_table = 23'b01110110000110110101101;
10'b1111000000: fsqrtinv_table = 23'b01110101111010010111010;
10'b1111000001: fsqrtinv_table = 23'b01110101101101111010010;
10'b1111000010: fsqrtinv_table = 23'b01110101100001011110011;
10'b1111000011: fsqrtinv_table = 23'b01110101010101000011111;
10'b1111000100: fsqrtinv_table = 23'b01110101001000101010100;
10'b1111000101: fsqrtinv_table = 23'b01110100111100010010011;
10'b1111000110: fsqrtinv_table = 23'b01110100101111111011100;
10'b1111000111: fsqrtinv_table = 23'b01110100100011100101111;
10'b1111001000: fsqrtinv_table = 23'b01110100010111010001100;
10'b1111001001: fsqrtinv_table = 23'b01110100001010111110010;
10'b1111001010: fsqrtinv_table = 23'b01110011111110101100010;
10'b1111001011: fsqrtinv_table = 23'b01110011110010011011100;
10'b1111001100: fsqrtinv_table = 23'b01110011100110001100000;
10'b1111001101: fsqrtinv_table = 23'b01110011011001111101101;
10'b1111001110: fsqrtinv_table = 23'b01110011001101110000100;
10'b1111001111: fsqrtinv_table = 23'b01110011000001100100100;
10'b1111010000: fsqrtinv_table = 23'b01110010110101011001110;
10'b1111010001: fsqrtinv_table = 23'b01110010101001010000010;
10'b1111010010: fsqrtinv_table = 23'b01110010011101000111111;
10'b1111010011: fsqrtinv_table = 23'b01110010010001000000110;
10'b1111010100: fsqrtinv_table = 23'b01110010000100111010110;
10'b1111010101: fsqrtinv_table = 23'b01110001111000110101111;
10'b1111010110: fsqrtinv_table = 23'b01110001101100110010011;
10'b1111010111: fsqrtinv_table = 23'b01110001100000101111111;
10'b1111011000: fsqrtinv_table = 23'b01110001010100101110101;
10'b1111011001: fsqrtinv_table = 23'b01110001001000101110100;
10'b1111011010: fsqrtinv_table = 23'b01110000111100101111101;
10'b1111011011: fsqrtinv_table = 23'b01110000110000110001111;
10'b1111011100: fsqrtinv_table = 23'b01110000100100110101010;
10'b1111011101: fsqrtinv_table = 23'b01110000011000111001111;
10'b1111011110: fsqrtinv_table = 23'b01110000001100111111101;
10'b1111011111: fsqrtinv_table = 23'b01110000000001000110100;
10'b1111100000: fsqrtinv_table = 23'b01101111110101001110100;
10'b1111100001: fsqrtinv_table = 23'b01101111101001010111101;
10'b1111100010: fsqrtinv_table = 23'b01101111011101100010000;
10'b1111100011: fsqrtinv_table = 23'b01101111010001101101100;
10'b1111100100: fsqrtinv_table = 23'b01101111000101111010000;
10'b1111100101: fsqrtinv_table = 23'b01101110111010000111110;
10'b1111100110: fsqrtinv_table = 23'b01101110101110010110101;
10'b1111100111: fsqrtinv_table = 23'b01101110100010100110101;
10'b1111101000: fsqrtinv_table = 23'b01101110010110110111111;
10'b1111101001: fsqrtinv_table = 23'b01101110001011001010001;
10'b1111101010: fsqrtinv_table = 23'b01101101111111011101100;
10'b1111101011: fsqrtinv_table = 23'b01101101110011110010000;
10'b1111101100: fsqrtinv_table = 23'b01101101101000000111101;
10'b1111101101: fsqrtinv_table = 23'b01101101011100011110011;
10'b1111101110: fsqrtinv_table = 23'b01101101010000110110001;
10'b1111101111: fsqrtinv_table = 23'b01101101000101001111001;
10'b1111110000: fsqrtinv_table = 23'b01101100111001101001010;
10'b1111110001: fsqrtinv_table = 23'b01101100101110000100011;
10'b1111110010: fsqrtinv_table = 23'b01101100100010100000101;
10'b1111110011: fsqrtinv_table = 23'b01101100010110111110000;
10'b1111110100: fsqrtinv_table = 23'b01101100001011011100100;
10'b1111110101: fsqrtinv_table = 23'b01101011111111111100000;
10'b1111110110: fsqrtinv_table = 23'b01101011110100011100101;
10'b1111110111: fsqrtinv_table = 23'b01101011101000111110011;
10'b1111111000: fsqrtinv_table = 23'b01101011011101100001001;
10'b1111111001: fsqrtinv_table = 23'b01101011010010000101001;
10'b1111111010: fsqrtinv_table = 23'b01101011000110101010000;
10'b1111111011: fsqrtinv_table = 23'b01101010111011010000001;
10'b1111111100: fsqrtinv_table = 23'b01101010101111110111010;
10'b1111111101: fsqrtinv_table = 23'b01101010100100011111011;
10'b1111111110: fsqrtinv_table = 23'b01101010011001001000101;
10'b1111111111: fsqrtinv_table = 23'b01101010001101110011000;

     endcase
    end
  endfunction

  wire [7:0] e1;
  wire [22:0] m1;
  assign e1 = x1[30:23];
  assign m1 = x1[22:0];

  wire [22:0] xs23, xsi23;
  assign xs23 = fsqrt_table({e1[0:0], m1[22:14]});
  assign xsi23 = fsqrtinv_table({e1[0:0], m1[22:14]});
  assign y1 = {1'b1, xs23};
  assign y2 = {1'b1, xsi23};

endmodule

`default_nettype wire
