`default_nettype none

module fdiv0(
  input wire [31:0] x2,
  output wire [23:0] y1,
  output wire [23:0] y2 );
  
  function [22:0] finv1 (
    input [11:0] m_input1 );
    begin
      case(m_input1)

12'b000000000000: finv1 = 23'b00000000000000000000000;
12'b000000000001: finv1 = 23'b11111111111000000000001;
12'b000000000010: finv1 = 23'b11111111110000000000100;
12'b000000000011: finv1 = 23'b11111111101000000001001;
12'b000000000100: finv1 = 23'b11111111100000000010000;
12'b000000000101: finv1 = 23'b11111111011000000011001;
12'b000000000110: finv1 = 23'b11111111010000000100100;
12'b000000000111: finv1 = 23'b11111111001000000110001;
12'b000000001000: finv1 = 23'b11111111000000001000000;
12'b000000001001: finv1 = 23'b11111110111000001010001;
12'b000000001010: finv1 = 23'b11111110110000001100100;
12'b000000001011: finv1 = 23'b11111110101000001111001;
12'b000000001100: finv1 = 23'b11111110100000010010000;
12'b000000001101: finv1 = 23'b11111110011000010101000;
12'b000000001110: finv1 = 23'b11111110010000011000011;
12'b000000001111: finv1 = 23'b11111110001000011100000;
12'b000000010000: finv1 = 23'b11111110000000011111111;
12'b000000010001: finv1 = 23'b11111101111000100100000;
12'b000000010010: finv1 = 23'b11111101110000101000011;
12'b000000010011: finv1 = 23'b11111101101000101100111;
12'b000000010100: finv1 = 23'b11111101100000110001110;
12'b000000010101: finv1 = 23'b11111101011000110110111;
12'b000000010110: finv1 = 23'b11111101010000111100001;
12'b000000010111: finv1 = 23'b11111101001001000001110;
12'b000000011000: finv1 = 23'b11111101000001000111101;
12'b000000011001: finv1 = 23'b11111100111001001101101;
12'b000000011010: finv1 = 23'b11111100110001010100000;
12'b000000011011: finv1 = 23'b11111100101001011010100;
12'b000000011100: finv1 = 23'b11111100100001100001011;
12'b000000011101: finv1 = 23'b11111100011001101000011;
12'b000000011110: finv1 = 23'b11111100010001101111101;
12'b000000011111: finv1 = 23'b11111100001001110111010;
12'b000000100000: finv1 = 23'b11111100000001111111000;
12'b000000100001: finv1 = 23'b11111011111010000111000;
12'b000000100010: finv1 = 23'b11111011110010001111010;
12'b000000100011: finv1 = 23'b11111011101010010111111;
12'b000000100100: finv1 = 23'b11111011100010100000101;
12'b000000100101: finv1 = 23'b11111011011010101001101;
12'b000000100110: finv1 = 23'b11111011010010110010111;
12'b000000100111: finv1 = 23'b11111011001010111100011;
12'b000000101000: finv1 = 23'b11111011000011000110001;
12'b000000101001: finv1 = 23'b11111010111011010000000;
12'b000000101010: finv1 = 23'b11111010110011011010010;
12'b000000101011: finv1 = 23'b11111010101011100100110;
12'b000000101100: finv1 = 23'b11111010100011101111011;
12'b000000101101: finv1 = 23'b11111010011011111010011;
12'b000000101110: finv1 = 23'b11111010010100000101101;
12'b000000101111: finv1 = 23'b11111010001100010001000;
12'b000000110000: finv1 = 23'b11111010000100011100101;
12'b000000110001: finv1 = 23'b11111001111100101000101;
12'b000000110010: finv1 = 23'b11111001110100110100110;
12'b000000110011: finv1 = 23'b11111001101101000001001;
12'b000000110100: finv1 = 23'b11111001100101001101110;
12'b000000110101: finv1 = 23'b11111001011101011010101;
12'b000000110110: finv1 = 23'b11111001010101100111110;
12'b000000110111: finv1 = 23'b11111001001101110101001;
12'b000000111000: finv1 = 23'b11111001000110000010110;
12'b000000111001: finv1 = 23'b11111000111110010000100;
12'b000000111010: finv1 = 23'b11111000110110011110101;
12'b000000111011: finv1 = 23'b11111000101110101101000;
12'b000000111100: finv1 = 23'b11111000100110111011100;
12'b000000111101: finv1 = 23'b11111000011111001010010;
12'b000000111110: finv1 = 23'b11111000010111011001011;
12'b000000111111: finv1 = 23'b11111000001111101000101;
12'b000001000000: finv1 = 23'b11111000000111111000001;
12'b000001000001: finv1 = 23'b11111000000000000111111;
12'b000001000010: finv1 = 23'b11110111111000010111111;
12'b000001000011: finv1 = 23'b11110111110000101000001;
12'b000001000100: finv1 = 23'b11110111101000111000100;
12'b000001000101: finv1 = 23'b11110111100001001001010;
12'b000001000110: finv1 = 23'b11110111011001011010010;
12'b000001000111: finv1 = 23'b11110111010001101011011;
12'b000001001000: finv1 = 23'b11110111001001111100110;
12'b000001001001: finv1 = 23'b11110111000010001110100;
12'b000001001010: finv1 = 23'b11110110111010100000011;
12'b000001001011: finv1 = 23'b11110110110010110010100;
12'b000001001100: finv1 = 23'b11110110101011000100111;
12'b000001001101: finv1 = 23'b11110110100011010111100;
12'b000001001110: finv1 = 23'b11110110011011101010010;
12'b000001001111: finv1 = 23'b11110110010011111101011;
12'b000001010000: finv1 = 23'b11110110001100010000101;
12'b000001010001: finv1 = 23'b11110110000100100100010;
12'b000001010010: finv1 = 23'b11110101111100111000000;
12'b000001010011: finv1 = 23'b11110101110101001100000;
12'b000001010100: finv1 = 23'b11110101101101100000010;
12'b000001010101: finv1 = 23'b11110101100101110100110;
12'b000001010110: finv1 = 23'b11110101011110001001100;
12'b000001010111: finv1 = 23'b11110101010110011110100;
12'b000001011000: finv1 = 23'b11110101001110110011101;
12'b000001011001: finv1 = 23'b11110101000111001001001;
12'b000001011010: finv1 = 23'b11110100111111011110110;
12'b000001011011: finv1 = 23'b11110100110111110100101;
12'b000001011100: finv1 = 23'b11110100110000001010110;
12'b000001011101: finv1 = 23'b11110100101000100001001;
12'b000001011110: finv1 = 23'b11110100100000110111110;
12'b000001011111: finv1 = 23'b11110100011001001110100;
12'b000001100000: finv1 = 23'b11110100010001100101101;
12'b000001100001: finv1 = 23'b11110100001001111100111;
12'b000001100010: finv1 = 23'b11110100000010010100100;
12'b000001100011: finv1 = 23'b11110011111010101100010;
12'b000001100100: finv1 = 23'b11110011110011000100010;
12'b000001100101: finv1 = 23'b11110011101011011100100;
12'b000001100110: finv1 = 23'b11110011100011110100111;
12'b000001100111: finv1 = 23'b11110011011100001101101;
12'b000001101000: finv1 = 23'b11110011010100100110100;
12'b000001101001: finv1 = 23'b11110011001100111111101;
12'b000001101010: finv1 = 23'b11110011000101011001001;
12'b000001101011: finv1 = 23'b11110010111101110010110;
12'b000001101100: finv1 = 23'b11110010110110001100100;
12'b000001101101: finv1 = 23'b11110010101110100110101;
12'b000001101110: finv1 = 23'b11110010100111000001000;
12'b000001101111: finv1 = 23'b11110010011111011011100;
12'b000001110000: finv1 = 23'b11110010010111110110010;
12'b000001110001: finv1 = 23'b11110010010000010001010;
12'b000001110010: finv1 = 23'b11110010001000101100100;
12'b000001110011: finv1 = 23'b11110010000001001000000;
12'b000001110100: finv1 = 23'b11110001111001100011101;
12'b000001110101: finv1 = 23'b11110001110001111111101;
12'b000001110110: finv1 = 23'b11110001101010011011110;
12'b000001110111: finv1 = 23'b11110001100010111000001;
12'b000001111000: finv1 = 23'b11110001011011010100110;
12'b000001111001: finv1 = 23'b11110001010011110001101;
12'b000001111010: finv1 = 23'b11110001001100001110110;
12'b000001111011: finv1 = 23'b11110001000100101100000;
12'b000001111100: finv1 = 23'b11110000111101001001100;
12'b000001111101: finv1 = 23'b11110000110101100111010;
12'b000001111110: finv1 = 23'b11110000101110000101010;
12'b000001111111: finv1 = 23'b11110000100110100011100;
12'b000010000000: finv1 = 23'b11110000011111000010000;
12'b000010000001: finv1 = 23'b11110000010111100000101;
12'b000010000010: finv1 = 23'b11110000001111111111100;
12'b000010000011: finv1 = 23'b11110000001000011110101;
12'b000010000100: finv1 = 23'b11110000000000111110000;
12'b000010000101: finv1 = 23'b11101111111001011101101;
12'b000010000110: finv1 = 23'b11101111110001111101011;
12'b000010000111: finv1 = 23'b11101111101010011101011;
12'b000010001000: finv1 = 23'b11101111100010111101110;
12'b000010001001: finv1 = 23'b11101111011011011110010;
12'b000010001010: finv1 = 23'b11101111010011111110111;
12'b000010001011: finv1 = 23'b11101111001100011111111;
12'b000010001100: finv1 = 23'b11101111000101000001000;
12'b000010001101: finv1 = 23'b11101110111101100010011;
12'b000010001110: finv1 = 23'b11101110110110000100000;
12'b000010001111: finv1 = 23'b11101110101110100101111;
12'b000010010000: finv1 = 23'b11101110100111001000000;
12'b000010010001: finv1 = 23'b11101110011111101010010;
12'b000010010010: finv1 = 23'b11101110011000001100110;
12'b000010010011: finv1 = 23'b11101110010000101111100;
12'b000010010100: finv1 = 23'b11101110001001010010100;
12'b000010010101: finv1 = 23'b11101110000001110101110;
12'b000010010110: finv1 = 23'b11101101111010011001001;
12'b000010010111: finv1 = 23'b11101101110010111100110;
12'b000010011000: finv1 = 23'b11101101101011100000101;
12'b000010011001: finv1 = 23'b11101101100100000100110;
12'b000010011010: finv1 = 23'b11101101011100101001001;
12'b000010011011: finv1 = 23'b11101101010101001101101;
12'b000010011100: finv1 = 23'b11101101001101110010011;
12'b000010011101: finv1 = 23'b11101101000110010111011;
12'b000010011110: finv1 = 23'b11101100111110111100101;
12'b000010011111: finv1 = 23'b11101100110111100010000;
12'b000010100000: finv1 = 23'b11101100110000000111110;
12'b000010100001: finv1 = 23'b11101100101000101101101;
12'b000010100010: finv1 = 23'b11101100100001010011110;
12'b000010100011: finv1 = 23'b11101100011001111010000;
12'b000010100100: finv1 = 23'b11101100010010100000101;
12'b000010100101: finv1 = 23'b11101100001011000111011;
12'b000010100110: finv1 = 23'b11101100000011101110011;
12'b000010100111: finv1 = 23'b11101011111100010101100;
12'b000010101000: finv1 = 23'b11101011110100111101000;
12'b000010101001: finv1 = 23'b11101011101101100100101;
12'b000010101010: finv1 = 23'b11101011100110001100100;
12'b000010101011: finv1 = 23'b11101011011110110100101;
12'b000010101100: finv1 = 23'b11101011010111011101000;
12'b000010101101: finv1 = 23'b11101011010000000101100;
12'b000010101110: finv1 = 23'b11101011001000101110010;
12'b000010101111: finv1 = 23'b11101011000001010111010;
12'b000010110000: finv1 = 23'b11101010111010000000100;
12'b000010110001: finv1 = 23'b11101010110010101001111;
12'b000010110010: finv1 = 23'b11101010101011010011100;
12'b000010110011: finv1 = 23'b11101010100011111101011;
12'b000010110100: finv1 = 23'b11101010011100100111100;
12'b000010110101: finv1 = 23'b11101010010101010001111;
12'b000010110110: finv1 = 23'b11101010001101111100011;
12'b000010110111: finv1 = 23'b11101010000110100111001;
12'b000010111000: finv1 = 23'b11101001111111010010001;
12'b000010111001: finv1 = 23'b11101001110111111101010;
12'b000010111010: finv1 = 23'b11101001110000101000101;
12'b000010111011: finv1 = 23'b11101001101001010100010;
12'b000010111100: finv1 = 23'b11101001100010000000001;
12'b000010111101: finv1 = 23'b11101001011010101100001;
12'b000010111110: finv1 = 23'b11101001010011011000100;
12'b000010111111: finv1 = 23'b11101001001100000101000;
12'b000011000000: finv1 = 23'b11101001000100110001101;
12'b000011000001: finv1 = 23'b11101000111101011110101;
12'b000011000010: finv1 = 23'b11101000110110001011110;
12'b000011000011: finv1 = 23'b11101000101110111001001;
12'b000011000100: finv1 = 23'b11101000100111100110110;
12'b000011000101: finv1 = 23'b11101000100000010100100;
12'b000011000110: finv1 = 23'b11101000011001000010100;
12'b000011000111: finv1 = 23'b11101000010001110000110;
12'b000011001000: finv1 = 23'b11101000001010011111010;
12'b000011001001: finv1 = 23'b11101000000011001101111;
12'b000011001010: finv1 = 23'b11100111111011111100110;
12'b000011001011: finv1 = 23'b11100111110100101011111;
12'b000011001100: finv1 = 23'b11100111101101011011010;
12'b000011001101: finv1 = 23'b11100111100110001010110;
12'b000011001110: finv1 = 23'b11100111011110111010100;
12'b000011001111: finv1 = 23'b11100111010111101010100;
12'b000011010000: finv1 = 23'b11100111010000011010101;
12'b000011010001: finv1 = 23'b11100111001001001011000;
12'b000011010010: finv1 = 23'b11100111000001111011101;
12'b000011010011: finv1 = 23'b11100110111010101100100;
12'b000011010100: finv1 = 23'b11100110110011011101100;
12'b000011010101: finv1 = 23'b11100110101100001110110;
12'b000011010110: finv1 = 23'b11100110100101000000010;
12'b000011010111: finv1 = 23'b11100110011101110010000;
12'b000011011000: finv1 = 23'b11100110010110100011111;
12'b000011011001: finv1 = 23'b11100110001111010110000;
12'b000011011010: finv1 = 23'b11100110001000001000010;
12'b000011011011: finv1 = 23'b11100110000000111010111;
12'b000011011100: finv1 = 23'b11100101111001101101101;
12'b000011011101: finv1 = 23'b11100101110010100000101;
12'b000011011110: finv1 = 23'b11100101101011010011110;
12'b000011011111: finv1 = 23'b11100101100100000111001;
12'b000011100000: finv1 = 23'b11100101011100111010110;
12'b000011100001: finv1 = 23'b11100101010101101110101;
12'b000011100010: finv1 = 23'b11100101001110100010101;
12'b000011100011: finv1 = 23'b11100101000111010110111;
12'b000011100100: finv1 = 23'b11100101000000001011011;
12'b000011100101: finv1 = 23'b11100100111001000000000;
12'b000011100110: finv1 = 23'b11100100110001110100111;
12'b000011100111: finv1 = 23'b11100100101010101010000;
12'b000011101000: finv1 = 23'b11100100100011011111011;
12'b000011101001: finv1 = 23'b11100100011100010100111;
12'b000011101010: finv1 = 23'b11100100010101001010101;
12'b000011101011: finv1 = 23'b11100100001110000000100;
12'b000011101100: finv1 = 23'b11100100000110110110110;
12'b000011101101: finv1 = 23'b11100011111111101101001;
12'b000011101110: finv1 = 23'b11100011111000100011101;
12'b000011101111: finv1 = 23'b11100011110001011010100;
12'b000011110000: finv1 = 23'b11100011101010010001100;
12'b000011110001: finv1 = 23'b11100011100011001000110;
12'b000011110010: finv1 = 23'b11100011011100000000001;
12'b000011110011: finv1 = 23'b11100011010100110111110;
12'b000011110100: finv1 = 23'b11100011001101101111101;
12'b000011110101: finv1 = 23'b11100011000110100111101;
12'b000011110110: finv1 = 23'b11100010111111011111111;
12'b000011110111: finv1 = 23'b11100010111000011000011;
12'b000011111000: finv1 = 23'b11100010110001010001001;
12'b000011111001: finv1 = 23'b11100010101010001010000;
12'b000011111010: finv1 = 23'b11100010100011000011001;
12'b000011111011: finv1 = 23'b11100010011011111100011;
12'b000011111100: finv1 = 23'b11100010010100110101111;
12'b000011111101: finv1 = 23'b11100010001101101111101;
12'b000011111110: finv1 = 23'b11100010000110101001101;
12'b000011111111: finv1 = 23'b11100001111111100011110;
12'b000100000000: finv1 = 23'b11100001111000011110001;
12'b000100000001: finv1 = 23'b11100001110001011000101;
12'b000100000010: finv1 = 23'b11100001101010010011100;
12'b000100000011: finv1 = 23'b11100001100011001110100;
12'b000100000100: finv1 = 23'b11100001011100001001101;
12'b000100000101: finv1 = 23'b11100001010101000101000;
12'b000100000110: finv1 = 23'b11100001001110000000101;
12'b000100000111: finv1 = 23'b11100001000110111100100;
12'b000100001000: finv1 = 23'b11100000111111111000100;
12'b000100001001: finv1 = 23'b11100000111000110100110;
12'b000100001010: finv1 = 23'b11100000110001110001001;
12'b000100001011: finv1 = 23'b11100000101010101101110;
12'b000100001100: finv1 = 23'b11100000100011101010101;
12'b000100001101: finv1 = 23'b11100000011100100111110;
12'b000100001110: finv1 = 23'b11100000010101100101000;
12'b000100001111: finv1 = 23'b11100000001110100010100;
12'b000100010000: finv1 = 23'b11100000000111100000001;
12'b000100010001: finv1 = 23'b11100000000000011110000;
12'b000100010010: finv1 = 23'b11011111111001011100001;
12'b000100010011: finv1 = 23'b11011111110010011010011;
12'b000100010100: finv1 = 23'b11011111101011011000111;
12'b000100010101: finv1 = 23'b11011111100100010111101;
12'b000100010110: finv1 = 23'b11011111011101010110100;
12'b000100010111: finv1 = 23'b11011111010110010101101;
12'b000100011000: finv1 = 23'b11011111001111010101000;
12'b000100011001: finv1 = 23'b11011111001000010100100;
12'b000100011010: finv1 = 23'b11011111000001010100010;
12'b000100011011: finv1 = 23'b11011110111010010100001;
12'b000100011100: finv1 = 23'b11011110110011010100010;
12'b000100011101: finv1 = 23'b11011110101100010100101;
12'b000100011110: finv1 = 23'b11011110100101010101001;
12'b000100011111: finv1 = 23'b11011110011110010101111;
12'b000100100000: finv1 = 23'b11011110010111010110111;
12'b000100100001: finv1 = 23'b11011110010000011000000;
12'b000100100010: finv1 = 23'b11011110001001011001011;
12'b000100100011: finv1 = 23'b11011110000010011011000;
12'b000100100100: finv1 = 23'b11011101111011011100110;
12'b000100100101: finv1 = 23'b11011101110100011110110;
12'b000100100110: finv1 = 23'b11011101101101100000111;
12'b000100100111: finv1 = 23'b11011101100110100011010;
12'b000100101000: finv1 = 23'b11011101011111100101111;
12'b000100101001: finv1 = 23'b11011101011000101000101;
12'b000100101010: finv1 = 23'b11011101010001101011101;
12'b000100101011: finv1 = 23'b11011101001010101110111;
12'b000100101100: finv1 = 23'b11011101000011110010010;
12'b000100101101: finv1 = 23'b11011100111100110101111;
12'b000100101110: finv1 = 23'b11011100110101111001101;
12'b000100101111: finv1 = 23'b11011100101110111101101;
12'b000100110000: finv1 = 23'b11011100101000000001111;
12'b000100110001: finv1 = 23'b11011100100001000110010;
12'b000100110010: finv1 = 23'b11011100011010001010111;
12'b000100110011: finv1 = 23'b11011100010011001111101;
12'b000100110100: finv1 = 23'b11011100001100010100110;
12'b000100110101: finv1 = 23'b11011100000101011001111;
12'b000100110110: finv1 = 23'b11011011111110011111011;
12'b000100110111: finv1 = 23'b11011011110111100100111;
12'b000100111000: finv1 = 23'b11011011110000101010110;
12'b000100111001: finv1 = 23'b11011011101001110000110;
12'b000100111010: finv1 = 23'b11011011100010110111000;
12'b000100111011: finv1 = 23'b11011011011011111101011;
12'b000100111100: finv1 = 23'b11011011010101000100000;
12'b000100111101: finv1 = 23'b11011011001110001010111;
12'b000100111110: finv1 = 23'b11011011000111010001111;
12'b000100111111: finv1 = 23'b11011011000000011001000;
12'b000101000000: finv1 = 23'b11011010111001100000100;
12'b000101000001: finv1 = 23'b11011010110010101000001;
12'b000101000010: finv1 = 23'b11011010101011101111111;
12'b000101000011: finv1 = 23'b11011010100100110111111;
12'b000101000100: finv1 = 23'b11011010011110000000001;
12'b000101000101: finv1 = 23'b11011010010111001000100;
12'b000101000110: finv1 = 23'b11011010010000010001001;
12'b000101000111: finv1 = 23'b11011010001001011010000;
12'b000101001000: finv1 = 23'b11011010000010100011000;
12'b000101001001: finv1 = 23'b11011001111011101100001;
12'b000101001010: finv1 = 23'b11011001110100110101100;
12'b000101001011: finv1 = 23'b11011001101101111111001;
12'b000101001100: finv1 = 23'b11011001100111001001000;
12'b000101001101: finv1 = 23'b11011001100000010011000;
12'b000101001110: finv1 = 23'b11011001011001011101001;
12'b000101001111: finv1 = 23'b11011001010010100111100;
12'b000101010000: finv1 = 23'b11011001001011110010001;
12'b000101010001: finv1 = 23'b11011001000100111100111;
12'b000101010010: finv1 = 23'b11011000111110000111111;
12'b000101010011: finv1 = 23'b11011000110111010011001;
12'b000101010100: finv1 = 23'b11011000110000011110100;
12'b000101010101: finv1 = 23'b11011000101001101010000;
12'b000101010110: finv1 = 23'b11011000100010110101111;
12'b000101010111: finv1 = 23'b11011000011100000001110;
12'b000101011000: finv1 = 23'b11011000010101001110000;
12'b000101011001: finv1 = 23'b11011000001110011010011;
12'b000101011010: finv1 = 23'b11011000000111100110111;
12'b000101011011: finv1 = 23'b11011000000000110011101;
12'b000101011100: finv1 = 23'b11010111111010000000101;
12'b000101011101: finv1 = 23'b11010111110011001101110;
12'b000101011110: finv1 = 23'b11010111101100011011001;
12'b000101011111: finv1 = 23'b11010111100101101000101;
12'b000101100000: finv1 = 23'b11010111011110110110011;
12'b000101100001: finv1 = 23'b11010111011000000100010;
12'b000101100010: finv1 = 23'b11010111010001010010011;
12'b000101100011: finv1 = 23'b11010111001010100000110;
12'b000101100100: finv1 = 23'b11010111000011101111010;
12'b000101100101: finv1 = 23'b11010110111100111101111;
12'b000101100110: finv1 = 23'b11010110110110001100111;
12'b000101100111: finv1 = 23'b11010110101111011011111;
12'b000101101000: finv1 = 23'b11010110101000101011010;
12'b000101101001: finv1 = 23'b11010110100001111010101;
12'b000101101010: finv1 = 23'b11010110011011001010011;
12'b000101101011: finv1 = 23'b11010110010100011010010;
12'b000101101100: finv1 = 23'b11010110001101101010010;
12'b000101101101: finv1 = 23'b11010110000110111010101;
12'b000101101110: finv1 = 23'b11010110000000001011000;
12'b000101101111: finv1 = 23'b11010101111001011011101;
12'b000101110000: finv1 = 23'b11010101110010101100100;
12'b000101110001: finv1 = 23'b11010101101011111101100;
12'b000101110010: finv1 = 23'b11010101100101001110110;
12'b000101110011: finv1 = 23'b11010101011110100000001;
12'b000101110100: finv1 = 23'b11010101010111110001110;
12'b000101110101: finv1 = 23'b11010101010001000011101;
12'b000101110110: finv1 = 23'b11010101001010010101101;
12'b000101110111: finv1 = 23'b11010101000011100111110;
12'b000101111000: finv1 = 23'b11010100111100111010001;
12'b000101111001: finv1 = 23'b11010100110110001100110;
12'b000101111010: finv1 = 23'b11010100101111011111100;
12'b000101111011: finv1 = 23'b11010100101000110010100;
12'b000101111100: finv1 = 23'b11010100100010000101101;
12'b000101111101: finv1 = 23'b11010100011011011001000;
12'b000101111110: finv1 = 23'b11010100010100101100100;
12'b000101111111: finv1 = 23'b11010100001110000000010;
12'b000110000000: finv1 = 23'b11010100000111010100001;
12'b000110000001: finv1 = 23'b11010100000000101000010;
12'b000110000010: finv1 = 23'b11010011111001111100100;
12'b000110000011: finv1 = 23'b11010011110011010001000;
12'b000110000100: finv1 = 23'b11010011101100100101101;
12'b000110000101: finv1 = 23'b11010011100101111010100;
12'b000110000110: finv1 = 23'b11010011011111001111101;
12'b000110000111: finv1 = 23'b11010011011000100100111;
12'b000110001000: finv1 = 23'b11010011010001111010010;
12'b000110001001: finv1 = 23'b11010011001011001111111;
12'b000110001010: finv1 = 23'b11010011000100100101110;
12'b000110001011: finv1 = 23'b11010010111101111011110;
12'b000110001100: finv1 = 23'b11010010110111010010000;
12'b000110001101: finv1 = 23'b11010010110000101000011;
12'b000110001110: finv1 = 23'b11010010101001111110111;
12'b000110001111: finv1 = 23'b11010010100011010101101;
12'b000110010000: finv1 = 23'b11010010011100101100101;
12'b000110010001: finv1 = 23'b11010010010110000011110;
12'b000110010010: finv1 = 23'b11010010001111011011001;
12'b000110010011: finv1 = 23'b11010010001000110010101;
12'b000110010100: finv1 = 23'b11010010000010001010011;
12'b000110010101: finv1 = 23'b11010001111011100010010;
12'b000110010110: finv1 = 23'b11010001110100111010011;
12'b000110010111: finv1 = 23'b11010001101110010010101;
12'b000110011000: finv1 = 23'b11010001100111101011001;
12'b000110011001: finv1 = 23'b11010001100001000011110;
12'b000110011010: finv1 = 23'b11010001011010011100101;
12'b000110011011: finv1 = 23'b11010001010011110101101;
12'b000110011100: finv1 = 23'b11010001001101001110111;
12'b000110011101: finv1 = 23'b11010001000110101000010;
12'b000110011110: finv1 = 23'b11010001000000000001111;
12'b000110011111: finv1 = 23'b11010000111001011011101;
12'b000110100000: finv1 = 23'b11010000110010110101100;
12'b000110100001: finv1 = 23'b11010000101100001111110;
12'b000110100010: finv1 = 23'b11010000100101101010000;
12'b000110100011: finv1 = 23'b11010000011111000100101;
12'b000110100100: finv1 = 23'b11010000011000011111010;
12'b000110100101: finv1 = 23'b11010000010001111010010;
12'b000110100110: finv1 = 23'b11010000001011010101010;
12'b000110100111: finv1 = 23'b11010000000100110000100;
12'b000110101000: finv1 = 23'b11001111111110001100000;
12'b000110101001: finv1 = 23'b11001111110111100111101;
12'b000110101010: finv1 = 23'b11001111110001000011100;
12'b000110101011: finv1 = 23'b11001111101010011111100;
12'b000110101100: finv1 = 23'b11001111100011111011110;
12'b000110101101: finv1 = 23'b11001111011101011000001;
12'b000110101110: finv1 = 23'b11001111010110110100101;
12'b000110101111: finv1 = 23'b11001111010000010001011;
12'b000110110000: finv1 = 23'b11001111001001101110011;
12'b000110110001: finv1 = 23'b11001111000011001011100;
12'b000110110010: finv1 = 23'b11001110111100101000110;
12'b000110110011: finv1 = 23'b11001110110110000110010;
12'b000110110100: finv1 = 23'b11001110101111100100000;
12'b000110110101: finv1 = 23'b11001110101001000001111;
12'b000110110110: finv1 = 23'b11001110100010011111111;
12'b000110110111: finv1 = 23'b11001110011011111110001;
12'b000110111000: finv1 = 23'b11001110010101011100100;
12'b000110111001: finv1 = 23'b11001110001110111011001;
12'b000110111010: finv1 = 23'b11001110001000011010000;
12'b000110111011: finv1 = 23'b11001110000001111000111;
12'b000110111100: finv1 = 23'b11001101111011011000001;
12'b000110111101: finv1 = 23'b11001101110100110111011;
12'b000110111110: finv1 = 23'b11001101101110010111000;
12'b000110111111: finv1 = 23'b11001101100111110110101;
12'b000111000000: finv1 = 23'b11001101100001010110100;
12'b000111000001: finv1 = 23'b11001101011010110110101;
12'b000111000010: finv1 = 23'b11001101010100010110111;
12'b000111000011: finv1 = 23'b11001101001101110111010;
12'b000111000100: finv1 = 23'b11001101000111010111111;
12'b000111000101: finv1 = 23'b11001101000000111000110;
12'b000111000110: finv1 = 23'b11001100111010011001110;
12'b000111000111: finv1 = 23'b11001100110011111010111;
12'b000111001000: finv1 = 23'b11001100101101011100010;
12'b000111001001: finv1 = 23'b11001100100110111101110;
12'b000111001010: finv1 = 23'b11001100100000011111100;
12'b000111001011: finv1 = 23'b11001100011010000001011;
12'b000111001100: finv1 = 23'b11001100010011100011100;
12'b000111001101: finv1 = 23'b11001100001101000101110;
12'b000111001110: finv1 = 23'b11001100000110101000001;
12'b000111001111: finv1 = 23'b11001100000000001010110;
12'b000111010000: finv1 = 23'b11001011111001101101101;
12'b000111010001: finv1 = 23'b11001011110011010000101;
12'b000111010010: finv1 = 23'b11001011101100110011110;
12'b000111010011: finv1 = 23'b11001011100110010111001;
12'b000111010100: finv1 = 23'b11001011011111111010101;
12'b000111010101: finv1 = 23'b11001011011001011110011;
12'b000111010110: finv1 = 23'b11001011010011000010010;
12'b000111010111: finv1 = 23'b11001011001100100110010;
12'b000111011000: finv1 = 23'b11001011000110001010100;
12'b000111011001: finv1 = 23'b11001010111111101111000;
12'b000111011010: finv1 = 23'b11001010111001010011101;
12'b000111011011: finv1 = 23'b11001010110010111000011;
12'b000111011100: finv1 = 23'b11001010101100011101011;
12'b000111011101: finv1 = 23'b11001010100110000010100;
12'b000111011110: finv1 = 23'b11001010011111100111111;
12'b000111011111: finv1 = 23'b11001010011001001101011;
12'b000111100000: finv1 = 23'b11001010010010110011000;
12'b000111100001: finv1 = 23'b11001010001100011000111;
12'b000111100010: finv1 = 23'b11001010000101111111000;
12'b000111100011: finv1 = 23'b11001001111111100101001;
12'b000111100100: finv1 = 23'b11001001111001001011101;
12'b000111100101: finv1 = 23'b11001001110010110010001;
12'b000111100110: finv1 = 23'b11001001101100011000111;
12'b000111100111: finv1 = 23'b11001001100101111111111;
12'b000111101000: finv1 = 23'b11001001011111100111000;
12'b000111101001: finv1 = 23'b11001001011001001110010;
12'b000111101010: finv1 = 23'b11001001010010110101110;
12'b000111101011: finv1 = 23'b11001001001100011101011;
12'b000111101100: finv1 = 23'b11001001000110000101010;
12'b000111101101: finv1 = 23'b11001000111111101101010;
12'b000111101110: finv1 = 23'b11001000111001010101100;
12'b000111101111: finv1 = 23'b11001000110010111101110;
12'b000111110000: finv1 = 23'b11001000101100100110011;
12'b000111110001: finv1 = 23'b11001000100110001111001;
12'b000111110010: finv1 = 23'b11001000011111111000000;
12'b000111110011: finv1 = 23'b11001000011001100001000;
12'b000111110100: finv1 = 23'b11001000010011001010010;
12'b000111110101: finv1 = 23'b11001000001100110011110;
12'b000111110110: finv1 = 23'b11001000000110011101011;
12'b000111110111: finv1 = 23'b11001000000000000111001;
12'b000111111000: finv1 = 23'b11000111111001110001001;
12'b000111111001: finv1 = 23'b11000111110011011011010;
12'b000111111010: finv1 = 23'b11000111101101000101100;
12'b000111111011: finv1 = 23'b11000111100110110000000;
12'b000111111100: finv1 = 23'b11000111100000011010110;
12'b000111111101: finv1 = 23'b11000111011010000101100;
12'b000111111110: finv1 = 23'b11000111010011110000100;
12'b000111111111: finv1 = 23'b11000111001101011011110;
12'b001000000000: finv1 = 23'b11000111000111000111001;
12'b001000000001: finv1 = 23'b11000111000000110010101;
12'b001000000010: finv1 = 23'b11000110111010011110011;
12'b001000000011: finv1 = 23'b11000110110100001010010;
12'b001000000100: finv1 = 23'b11000110101101110110011;
12'b001000000101: finv1 = 23'b11000110100111100010101;
12'b001000000110: finv1 = 23'b11000110100001001111000;
12'b001000000111: finv1 = 23'b11000110011010111011101;
12'b001000001000: finv1 = 23'b11000110010100101000011;
12'b001000001001: finv1 = 23'b11000110001110010101011;
12'b001000001010: finv1 = 23'b11000110001000000010100;
12'b001000001011: finv1 = 23'b11000110000001101111110;
12'b001000001100: finv1 = 23'b11000101111011011101010;
12'b001000001101: finv1 = 23'b11000101110101001010111;
12'b001000001110: finv1 = 23'b11000101101110111000101;
12'b001000001111: finv1 = 23'b11000101101000100110101;
12'b001000010000: finv1 = 23'b11000101100010010100111;
12'b001000010001: finv1 = 23'b11000101011100000011001;
12'b001000010010: finv1 = 23'b11000101010101110001101;
12'b001000010011: finv1 = 23'b11000101001111100000011;
12'b001000010100: finv1 = 23'b11000101001001001111010;
12'b001000010101: finv1 = 23'b11000101000010111110010;
12'b001000010110: finv1 = 23'b11000100111100101101100;
12'b001000010111: finv1 = 23'b11000100110110011100111;
12'b001000011000: finv1 = 23'b11000100110000001100011;
12'b001000011001: finv1 = 23'b11000100101001111100001;
12'b001000011010: finv1 = 23'b11000100100011101100000;
12'b001000011011: finv1 = 23'b11000100011101011100001;
12'b001000011100: finv1 = 23'b11000100010111001100011;
12'b001000011101: finv1 = 23'b11000100010000111100110;
12'b001000011110: finv1 = 23'b11000100001010101101011;
12'b001000011111: finv1 = 23'b11000100000100011110001;
12'b001000100000: finv1 = 23'b11000011111110001111000;
12'b001000100001: finv1 = 23'b11000011111000000000001;
12'b001000100010: finv1 = 23'b11000011110001110001011;
12'b001000100011: finv1 = 23'b11000011101011100010111;
12'b001000100100: finv1 = 23'b11000011100101010100100;
12'b001000100101: finv1 = 23'b11000011011111000110010;
12'b001000100110: finv1 = 23'b11000011011000111000010;
12'b001000100111: finv1 = 23'b11000011010010101010011;
12'b001000101000: finv1 = 23'b11000011001100011100101;
12'b001000101001: finv1 = 23'b11000011000110001111001;
12'b001000101010: finv1 = 23'b11000011000000000001110;
12'b001000101011: finv1 = 23'b11000010111001110100101;
12'b001000101100: finv1 = 23'b11000010110011100111101;
12'b001000101101: finv1 = 23'b11000010101101011010110;
12'b001000101110: finv1 = 23'b11000010100111001110000;
12'b001000101111: finv1 = 23'b11000010100001000001100;
12'b001000110000: finv1 = 23'b11000010011010110101010;
12'b001000110001: finv1 = 23'b11000010010100101001001;
12'b001000110010: finv1 = 23'b11000010001110011101001;
12'b001000110011: finv1 = 23'b11000010001000010001010;
12'b001000110100: finv1 = 23'b11000010000010000101101;
12'b001000110101: finv1 = 23'b11000001111011111010001;
12'b001000110110: finv1 = 23'b11000001110101101110111;
12'b001000110111: finv1 = 23'b11000001101111100011101;
12'b001000111000: finv1 = 23'b11000001101001011000110;
12'b001000111001: finv1 = 23'b11000001100011001101111;
12'b001000111010: finv1 = 23'b11000001011101000011010;
12'b001000111011: finv1 = 23'b11000001010110111000110;
12'b001000111100: finv1 = 23'b11000001010000101110100;
12'b001000111101: finv1 = 23'b11000001001010100100011;
12'b001000111110: finv1 = 23'b11000001000100011010011;
12'b001000111111: finv1 = 23'b11000000111110010000101;
12'b001001000000: finv1 = 23'b11000000111000000111000;
12'b001001000001: finv1 = 23'b11000000110001111101100;
12'b001001000010: finv1 = 23'b11000000101011110100010;
12'b001001000011: finv1 = 23'b11000000100101101011001;
12'b001001000100: finv1 = 23'b11000000011111100010010;
12'b001001000101: finv1 = 23'b11000000011001011001100;
12'b001001000110: finv1 = 23'b11000000010011010000111;
12'b001001000111: finv1 = 23'b11000000001101001000011;
12'b001001001000: finv1 = 23'b11000000000111000000001;
12'b001001001001: finv1 = 23'b11000000000000111000000;
12'b001001001010: finv1 = 23'b10111111111010110000000;
12'b001001001011: finv1 = 23'b10111111110100101000010;
12'b001001001100: finv1 = 23'b10111111101110100000101;
12'b001001001101: finv1 = 23'b10111111101000011001010;
12'b001001001110: finv1 = 23'b10111111100010010010000;
12'b001001001111: finv1 = 23'b10111111011100001010111;
12'b001001010000: finv1 = 23'b10111111010110000011111;
12'b001001010001: finv1 = 23'b10111111001111111101001;
12'b001001010010: finv1 = 23'b10111111001001110110100;
12'b001001010011: finv1 = 23'b10111111000011110000001;
12'b001001010100: finv1 = 23'b10111110111101101001111;
12'b001001010101: finv1 = 23'b10111110110111100011110;
12'b001001010110: finv1 = 23'b10111110110001011101110;
12'b001001010111: finv1 = 23'b10111110101011011000000;
12'b001001011000: finv1 = 23'b10111110100101010010011;
12'b001001011001: finv1 = 23'b10111110011111001101000;
12'b001001011010: finv1 = 23'b10111110011001000111110;
12'b001001011011: finv1 = 23'b10111110010011000010101;
12'b001001011100: finv1 = 23'b10111110001100111101101;
12'b001001011101: finv1 = 23'b10111110000110111000111;
12'b001001011110: finv1 = 23'b10111110000000110100010;
12'b001001011111: finv1 = 23'b10111101111010101111111;
12'b001001100000: finv1 = 23'b10111101110100101011100;
12'b001001100001: finv1 = 23'b10111101101110100111011;
12'b001001100010: finv1 = 23'b10111101101000100011100;
12'b001001100011: finv1 = 23'b10111101100010011111101;
12'b001001100100: finv1 = 23'b10111101011100011100000;
12'b001001100101: finv1 = 23'b10111101010110011000101;
12'b001001100110: finv1 = 23'b10111101010000010101010;
12'b001001100111: finv1 = 23'b10111101001010010010001;
12'b001001101000: finv1 = 23'b10111101000100001111010;
12'b001001101001: finv1 = 23'b10111100111110001100011;
12'b001001101010: finv1 = 23'b10111100111000001001110;
12'b001001101011: finv1 = 23'b10111100110010000111010;
12'b001001101100: finv1 = 23'b10111100101100000101000;
12'b001001101101: finv1 = 23'b10111100100110000010111;
12'b001001101110: finv1 = 23'b10111100100000000000111;
12'b001001101111: finv1 = 23'b10111100011001111111000;
12'b001001110000: finv1 = 23'b10111100010011111101011;
12'b001001110001: finv1 = 23'b10111100001101111011111;
12'b001001110010: finv1 = 23'b10111100000111111010101;
12'b001001110011: finv1 = 23'b10111100000001111001011;
12'b001001110100: finv1 = 23'b10111011111011111000011;
12'b001001110101: finv1 = 23'b10111011110101110111101;
12'b001001110110: finv1 = 23'b10111011101111110110111;
12'b001001110111: finv1 = 23'b10111011101001110110011;
12'b001001111000: finv1 = 23'b10111011100011110110000;
12'b001001111001: finv1 = 23'b10111011011101110101111;
12'b001001111010: finv1 = 23'b10111011010111110101111;
12'b001001111011: finv1 = 23'b10111011010001110110000;
12'b001001111100: finv1 = 23'b10111011001011110110010;
12'b001001111101: finv1 = 23'b10111011000101110110110;
12'b001001111110: finv1 = 23'b10111010111111110111011;
12'b001001111111: finv1 = 23'b10111010111001111000001;
12'b001010000000: finv1 = 23'b10111010110011111001001;
12'b001010000001: finv1 = 23'b10111010101101111010010;
12'b001010000010: finv1 = 23'b10111010100111111011100;
12'b001010000011: finv1 = 23'b10111010100001111100111;
12'b001010000100: finv1 = 23'b10111010011011111110100;
12'b001010000101: finv1 = 23'b10111010010110000000010;
12'b001010000110: finv1 = 23'b10111010010000000010001;
12'b001010000111: finv1 = 23'b10111010001010000100010;
12'b001010001000: finv1 = 23'b10111010000100000110100;
12'b001010001001: finv1 = 23'b10111001111110001000111;
12'b001010001010: finv1 = 23'b10111001111000001011011;
12'b001010001011: finv1 = 23'b10111001110010001110001;
12'b001010001100: finv1 = 23'b10111001101100010001000;
12'b001010001101: finv1 = 23'b10111001100110010100001;
12'b001010001110: finv1 = 23'b10111001100000010111010;
12'b001010001111: finv1 = 23'b10111001011010011010101;
12'b001010010000: finv1 = 23'b10111001010100011110001;
12'b001010010001: finv1 = 23'b10111001001110100001111;
12'b001010010010: finv1 = 23'b10111001001000100101110;
12'b001010010011: finv1 = 23'b10111001000010101001110;
12'b001010010100: finv1 = 23'b10111000111100101101111;
12'b001010010101: finv1 = 23'b10111000110110110010001;
12'b001010010110: finv1 = 23'b10111000110000110110101;
12'b001010010111: finv1 = 23'b10111000101010111011010;
12'b001010011000: finv1 = 23'b10111000100101000000001;
12'b001010011001: finv1 = 23'b10111000011111000101001;
12'b001010011010: finv1 = 23'b10111000011001001010001;
12'b001010011011: finv1 = 23'b10111000010011001111100;
12'b001010011100: finv1 = 23'b10111000001101010100111;
12'b001010011101: finv1 = 23'b10111000000111011010100;
12'b001010011110: finv1 = 23'b10111000000001100000010;
12'b001010011111: finv1 = 23'b10110111111011100110001;
12'b001010100000: finv1 = 23'b10110111110101101100010;
12'b001010100001: finv1 = 23'b10110111101111110010100;
12'b001010100010: finv1 = 23'b10110111101001111000111;
12'b001010100011: finv1 = 23'b10110111100011111111011;
12'b001010100100: finv1 = 23'b10110111011110000110001;
12'b001010100101: finv1 = 23'b10110111011000001101000;
12'b001010100110: finv1 = 23'b10110111010010010100000;
12'b001010100111: finv1 = 23'b10110111001100011011001;
12'b001010101000: finv1 = 23'b10110111000110100010100;
12'b001010101001: finv1 = 23'b10110111000000101010000;
12'b001010101010: finv1 = 23'b10110110111010110001101;
12'b001010101011: finv1 = 23'b10110110110100111001100;
12'b001010101100: finv1 = 23'b10110110101111000001100;
12'b001010101101: finv1 = 23'b10110110101001001001101;
12'b001010101110: finv1 = 23'b10110110100011010001111;
12'b001010101111: finv1 = 23'b10110110011101011010010;
12'b001010110000: finv1 = 23'b10110110010111100010111;
12'b001010110001: finv1 = 23'b10110110010001101011101;
12'b001010110010: finv1 = 23'b10110110001011110100100;
12'b001010110011: finv1 = 23'b10110110000101111101101;
12'b001010110100: finv1 = 23'b10110110000000000110111;
12'b001010110101: finv1 = 23'b10110101111010010000010;
12'b001010110110: finv1 = 23'b10110101110100011001110;
12'b001010110111: finv1 = 23'b10110101101110100011100;
12'b001010111000: finv1 = 23'b10110101101000101101010;
12'b001010111001: finv1 = 23'b10110101100010110111010;
12'b001010111010: finv1 = 23'b10110101011101000001100;
12'b001010111011: finv1 = 23'b10110101010111001011110;
12'b001010111100: finv1 = 23'b10110101010001010110010;
12'b001010111101: finv1 = 23'b10110101001011100000111;
12'b001010111110: finv1 = 23'b10110101000101101011101;
12'b001010111111: finv1 = 23'b10110100111111110110101;
12'b001011000000: finv1 = 23'b10110100111010000001110;
12'b001011000001: finv1 = 23'b10110100110100001101000;
12'b001011000010: finv1 = 23'b10110100101110011000011;
12'b001011000011: finv1 = 23'b10110100101000100011111;
12'b001011000100: finv1 = 23'b10110100100010101111101;
12'b001011000101: finv1 = 23'b10110100011100111011100;
12'b001011000110: finv1 = 23'b10110100010111000111100;
12'b001011000111: finv1 = 23'b10110100010001010011110;
12'b001011001000: finv1 = 23'b10110100001011100000000;
12'b001011001001: finv1 = 23'b10110100000101101100100;
12'b001011001010: finv1 = 23'b10110011111111111001010;
12'b001011001011: finv1 = 23'b10110011111010000110000;
12'b001011001100: finv1 = 23'b10110011110100010011000;
12'b001011001101: finv1 = 23'b10110011101110100000000;
12'b001011001110: finv1 = 23'b10110011101000101101010;
12'b001011001111: finv1 = 23'b10110011100010111010110;
12'b001011010000: finv1 = 23'b10110011011101001000010;
12'b001011010001: finv1 = 23'b10110011010111010110000;
12'b001011010010: finv1 = 23'b10110011010001100011111;
12'b001011010011: finv1 = 23'b10110011001011110001111;
12'b001011010100: finv1 = 23'b10110011000110000000001;
12'b001011010101: finv1 = 23'b10110011000000001110100;
12'b001011010110: finv1 = 23'b10110010111010011100111;
12'b001011010111: finv1 = 23'b10110010110100101011101;
12'b001011011000: finv1 = 23'b10110010101110111010011;
12'b001011011001: finv1 = 23'b10110010101001001001011;
12'b001011011010: finv1 = 23'b10110010100011011000011;
12'b001011011011: finv1 = 23'b10110010011101100111101;
12'b001011011100: finv1 = 23'b10110010010111110111001;
12'b001011011101: finv1 = 23'b10110010010010000110101;
12'b001011011110: finv1 = 23'b10110010001100010110011;
12'b001011011111: finv1 = 23'b10110010000110100110010;
12'b001011100000: finv1 = 23'b10110010000000110110010;
12'b001011100001: finv1 = 23'b10110001111011000110011;
12'b001011100010: finv1 = 23'b10110001110101010110110;
12'b001011100011: finv1 = 23'b10110001101111100111010;
12'b001011100100: finv1 = 23'b10110001101001110111111;
12'b001011100101: finv1 = 23'b10110001100100001000101;
12'b001011100110: finv1 = 23'b10110001011110011001100;
12'b001011100111: finv1 = 23'b10110001011000101010101;
12'b001011101000: finv1 = 23'b10110001010010111011111;
12'b001011101001: finv1 = 23'b10110001001101001101010;
12'b001011101010: finv1 = 23'b10110001000111011110110;
12'b001011101011: finv1 = 23'b10110001000001110000100;
12'b001011101100: finv1 = 23'b10110000111100000010011;
12'b001011101101: finv1 = 23'b10110000110110010100011;
12'b001011101110: finv1 = 23'b10110000110000100110100;
12'b001011101111: finv1 = 23'b10110000101010111000110;
12'b001011110000: finv1 = 23'b10110000100101001011010;
12'b001011110001: finv1 = 23'b10110000011111011101110;
12'b001011110010: finv1 = 23'b10110000011001110000100;
12'b001011110011: finv1 = 23'b10110000010100000011011;
12'b001011110100: finv1 = 23'b10110000001110010110100;
12'b001011110101: finv1 = 23'b10110000001000101001101;
12'b001011110110: finv1 = 23'b10110000000010111101000;
12'b001011110111: finv1 = 23'b10101111111101010000100;
12'b001011111000: finv1 = 23'b10101111110111100100001;
12'b001011111001: finv1 = 23'b10101111110001111000000;
12'b001011111010: finv1 = 23'b10101111101100001011111;
12'b001011111011: finv1 = 23'b10101111100110100000000;
12'b001011111100: finv1 = 23'b10101111100000110100010;
12'b001011111101: finv1 = 23'b10101111011011001000101;
12'b001011111110: finv1 = 23'b10101111010101011101010;
12'b001011111111: finv1 = 23'b10101111001111110001111;
12'b001100000000: finv1 = 23'b10101111001010000110110;
12'b001100000001: finv1 = 23'b10101111000100011011110;
12'b001100000010: finv1 = 23'b10101110111110110000111;
12'b001100000011: finv1 = 23'b10101110111001000110001;
12'b001100000100: finv1 = 23'b10101110110011011011101;
12'b001100000101: finv1 = 23'b10101110101101110001010;
12'b001100000110: finv1 = 23'b10101110101000000111000;
12'b001100000111: finv1 = 23'b10101110100010011100111;
12'b001100001000: finv1 = 23'b10101110011100110010111;
12'b001100001001: finv1 = 23'b10101110010111001001000;
12'b001100001010: finv1 = 23'b10101110010001011111011;
12'b001100001011: finv1 = 23'b10101110001011110101111;
12'b001100001100: finv1 = 23'b10101110000110001100100;
12'b001100001101: finv1 = 23'b10101110000000100011010;
12'b001100001110: finv1 = 23'b10101101111010111010010;
12'b001100001111: finv1 = 23'b10101101110101010001010;
12'b001100010000: finv1 = 23'b10101101101111101000100;
12'b001100010001: finv1 = 23'b10101101101001111111111;
12'b001100010010: finv1 = 23'b10101101100100010111011;
12'b001100010011: finv1 = 23'b10101101011110101111000;
12'b001100010100: finv1 = 23'b10101101011001000110111;
12'b001100010101: finv1 = 23'b10101101010011011110111;
12'b001100010110: finv1 = 23'b10101101001101110110111;
12'b001100010111: finv1 = 23'b10101101001000001111010;
12'b001100011000: finv1 = 23'b10101101000010100111101;
12'b001100011001: finv1 = 23'b10101100111101000000001;
12'b001100011010: finv1 = 23'b10101100110111011000111;
12'b001100011011: finv1 = 23'b10101100110001110001101;
12'b001100011100: finv1 = 23'b10101100101100001010101;
12'b001100011101: finv1 = 23'b10101100100110100011111;
12'b001100011110: finv1 = 23'b10101100100000111101001;
12'b001100011111: finv1 = 23'b10101100011011010110100;
12'b001100100000: finv1 = 23'b10101100010101110000001;
12'b001100100001: finv1 = 23'b10101100010000001001111;
12'b001100100010: finv1 = 23'b10101100001010100011110;
12'b001100100011: finv1 = 23'b10101100000100111101110;
12'b001100100100: finv1 = 23'b10101011111111010111111;
12'b001100100101: finv1 = 23'b10101011111001110010001;
12'b001100100110: finv1 = 23'b10101011110100001100101;
12'b001100100111: finv1 = 23'b10101011101110100111010;
12'b001100101000: finv1 = 23'b10101011101001000010000;
12'b001100101001: finv1 = 23'b10101011100011011100111;
12'b001100101010: finv1 = 23'b10101011011101110111111;
12'b001100101011: finv1 = 23'b10101011011000010011001;
12'b001100101100: finv1 = 23'b10101011010010101110011;
12'b001100101101: finv1 = 23'b10101011001101001001111;
12'b001100101110: finv1 = 23'b10101011000111100101100;
12'b001100101111: finv1 = 23'b10101011000010000001010;
12'b001100110000: finv1 = 23'b10101010111100011101001;
12'b001100110001: finv1 = 23'b10101010110110111001010;
12'b001100110010: finv1 = 23'b10101010110001010101100;
12'b001100110011: finv1 = 23'b10101010101011110001110;
12'b001100110100: finv1 = 23'b10101010100110001110010;
12'b001100110101: finv1 = 23'b10101010100000101010111;
12'b001100110110: finv1 = 23'b10101010011011000111101;
12'b001100110111: finv1 = 23'b10101010010101100100101;
12'b001100111000: finv1 = 23'b10101010010000000001101;
12'b001100111001: finv1 = 23'b10101010001010011110111;
12'b001100111010: finv1 = 23'b10101010000100111100010;
12'b001100111011: finv1 = 23'b10101001111111011001110;
12'b001100111100: finv1 = 23'b10101001111001110111011;
12'b001100111101: finv1 = 23'b10101001110100010101001;
12'b001100111110: finv1 = 23'b10101001101110110011001;
12'b001100111111: finv1 = 23'b10101001101001010001001;
12'b001101000000: finv1 = 23'b10101001100011101111011;
12'b001101000001: finv1 = 23'b10101001011110001101110;
12'b001101000010: finv1 = 23'b10101001011000101100010;
12'b001101000011: finv1 = 23'b10101001010011001010111;
12'b001101000100: finv1 = 23'b10101001001101101001101;
12'b001101000101: finv1 = 23'b10101001001000001000101;
12'b001101000110: finv1 = 23'b10101001000010100111110;
12'b001101000111: finv1 = 23'b10101000111101000110111;
12'b001101001000: finv1 = 23'b10101000110111100110010;
12'b001101001001: finv1 = 23'b10101000110010000101110;
12'b001101001010: finv1 = 23'b10101000101100100101011;
12'b001101001011: finv1 = 23'b10101000100111000101010;
12'b001101001100: finv1 = 23'b10101000100001100101001;
12'b001101001101: finv1 = 23'b10101000011100000101010;
12'b001101001110: finv1 = 23'b10101000010110100101100;
12'b001101001111: finv1 = 23'b10101000010001000101111;
12'b001101010000: finv1 = 23'b10101000001011100110011;
12'b001101010001: finv1 = 23'b10101000000110000111000;
12'b001101010010: finv1 = 23'b10101000000000100111110;
12'b001101010011: finv1 = 23'b10100111111011001000101;
12'b001101010100: finv1 = 23'b10100111110101101001110;
12'b001101010101: finv1 = 23'b10100111110000001011000;
12'b001101010110: finv1 = 23'b10100111101010101100011;
12'b001101010111: finv1 = 23'b10100111100101001101111;
12'b001101011000: finv1 = 23'b10100111011111101111100;
12'b001101011001: finv1 = 23'b10100111011010010001010;
12'b001101011010: finv1 = 23'b10100111010100110011001;
12'b001101011011: finv1 = 23'b10100111001111010101010;
12'b001101011100: finv1 = 23'b10100111001001110111011;
12'b001101011101: finv1 = 23'b10100111000100011001110;
12'b001101011110: finv1 = 23'b10100110111110111100010;
12'b001101011111: finv1 = 23'b10100110111001011110111;
12'b001101100000: finv1 = 23'b10100110110100000001101;
12'b001101100001: finv1 = 23'b10100110101110100100100;
12'b001101100010: finv1 = 23'b10100110101001000111101;
12'b001101100011: finv1 = 23'b10100110100011101010110;
12'b001101100100: finv1 = 23'b10100110011110001110001;
12'b001101100101: finv1 = 23'b10100110011000110001101;
12'b001101100110: finv1 = 23'b10100110010011010101010;
12'b001101100111: finv1 = 23'b10100110001101111001000;
12'b001101101000: finv1 = 23'b10100110001000011100111;
12'b001101101001: finv1 = 23'b10100110000011000000111;
12'b001101101010: finv1 = 23'b10100101111101100101000;
12'b001101101011: finv1 = 23'b10100101111000001001011;
12'b001101101100: finv1 = 23'b10100101110010101101111;
12'b001101101101: finv1 = 23'b10100101101101010010011;
12'b001101101110: finv1 = 23'b10100101100111110111001;
12'b001101101111: finv1 = 23'b10100101100010011100000;
12'b001101110000: finv1 = 23'b10100101011101000001000;
12'b001101110001: finv1 = 23'b10100101010111100110001;
12'b001101110010: finv1 = 23'b10100101010010001011100;
12'b001101110011: finv1 = 23'b10100101001100110000111;
12'b001101110100: finv1 = 23'b10100101000111010110100;
12'b001101110101: finv1 = 23'b10100101000001111100001;
12'b001101110110: finv1 = 23'b10100100111100100010000;
12'b001101110111: finv1 = 23'b10100100110111001000000;
12'b001101111000: finv1 = 23'b10100100110001101110001;
12'b001101111001: finv1 = 23'b10100100101100010100011;
12'b001101111010: finv1 = 23'b10100100100110111010110;
12'b001101111011: finv1 = 23'b10100100100001100001011;
12'b001101111100: finv1 = 23'b10100100011100001000000;
12'b001101111101: finv1 = 23'b10100100010110101110111;
12'b001101111110: finv1 = 23'b10100100010001010101110;
12'b001101111111: finv1 = 23'b10100100001011111100111;
12'b001110000000: finv1 = 23'b10100100000110100100001;
12'b001110000001: finv1 = 23'b10100100000001001011100;
12'b001110000010: finv1 = 23'b10100011111011110011000;
12'b001110000011: finv1 = 23'b10100011110110011010101;
12'b001110000100: finv1 = 23'b10100011110001000010011;
12'b001110000101: finv1 = 23'b10100011101011101010011;
12'b001110000110: finv1 = 23'b10100011100110010010011;
12'b001110000111: finv1 = 23'b10100011100000111010101;
12'b001110001000: finv1 = 23'b10100011011011100010111;
12'b001110001001: finv1 = 23'b10100011010110001011011;
12'b001110001010: finv1 = 23'b10100011010000110100000;
12'b001110001011: finv1 = 23'b10100011001011011100110;
12'b001110001100: finv1 = 23'b10100011000110000101101;
12'b001110001101: finv1 = 23'b10100011000000101110101;
12'b001110001110: finv1 = 23'b10100010111011010111110;
12'b001110001111: finv1 = 23'b10100010110110000001001;
12'b001110010000: finv1 = 23'b10100010110000101010100;
12'b001110010001: finv1 = 23'b10100010101011010100001;
12'b001110010010: finv1 = 23'b10100010100101111101110;
12'b001110010011: finv1 = 23'b10100010100000100111101;
12'b001110010100: finv1 = 23'b10100010011011010001101;
12'b001110010101: finv1 = 23'b10100010010101111011110;
12'b001110010110: finv1 = 23'b10100010010000100110000;
12'b001110010111: finv1 = 23'b10100010001011010000011;
12'b001110011000: finv1 = 23'b10100010000101111010111;
12'b001110011001: finv1 = 23'b10100010000000100101100;
12'b001110011010: finv1 = 23'b10100001111011010000011;
12'b001110011011: finv1 = 23'b10100001110101111011010;
12'b001110011100: finv1 = 23'b10100001110000100110011;
12'b001110011101: finv1 = 23'b10100001101011010001100;
12'b001110011110: finv1 = 23'b10100001100101111100111;
12'b001110011111: finv1 = 23'b10100001100000101000011;
12'b001110100000: finv1 = 23'b10100001011011010100000;
12'b001110100001: finv1 = 23'b10100001010101111111110;
12'b001110100010: finv1 = 23'b10100001010000101011101;
12'b001110100011: finv1 = 23'b10100001001011010111101;
12'b001110100100: finv1 = 23'b10100001000110000011110;
12'b001110100101: finv1 = 23'b10100001000000110000000;
12'b001110100110: finv1 = 23'b10100000111011011100100;
12'b001110100111: finv1 = 23'b10100000110110001001000;
12'b001110101000: finv1 = 23'b10100000110000110101110;
12'b001110101001: finv1 = 23'b10100000101011100010100;
12'b001110101010: finv1 = 23'b10100000100110001111100;
12'b001110101011: finv1 = 23'b10100000100000111100101;
12'b001110101100: finv1 = 23'b10100000011011101001111;
12'b001110101101: finv1 = 23'b10100000010110010111010;
12'b001110101110: finv1 = 23'b10100000010001000100110;
12'b001110101111: finv1 = 23'b10100000001011110010011;
12'b001110110000: finv1 = 23'b10100000000110100000001;
12'b001110110001: finv1 = 23'b10100000000001001110000;
12'b001110110010: finv1 = 23'b10011111111011111100000;
12'b001110110011: finv1 = 23'b10011111110110101010010;
12'b001110110100: finv1 = 23'b10011111110001011000100;
12'b001110110101: finv1 = 23'b10011111101100000111000;
12'b001110110110: finv1 = 23'b10011111100110110101100;
12'b001110110111: finv1 = 23'b10011111100001100100010;
12'b001110111000: finv1 = 23'b10011111011100010011001;
12'b001110111001: finv1 = 23'b10011111010111000010000;
12'b001110111010: finv1 = 23'b10011111010001110001001;
12'b001110111011: finv1 = 23'b10011111001100100000011;
12'b001110111100: finv1 = 23'b10011111000111001111110;
12'b001110111101: finv1 = 23'b10011111000001111111010;
12'b001110111110: finv1 = 23'b10011110111100101110111;
12'b001110111111: finv1 = 23'b10011110110111011110101;
12'b001111000000: finv1 = 23'b10011110110010001110101;
12'b001111000001: finv1 = 23'b10011110101100111110101;
12'b001111000010: finv1 = 23'b10011110100111101110110;
12'b001111000011: finv1 = 23'b10011110100010011111001;
12'b001111000100: finv1 = 23'b10011110011101001111100;
12'b001111000101: finv1 = 23'b10011110011000000000001;
12'b001111000110: finv1 = 23'b10011110010010110000110;
12'b001111000111: finv1 = 23'b10011110001101100001101;
12'b001111001000: finv1 = 23'b10011110001000010010101;
12'b001111001001: finv1 = 23'b10011110000011000011110;
12'b001111001010: finv1 = 23'b10011101111101110100111;
12'b001111001011: finv1 = 23'b10011101111000100110010;
12'b001111001100: finv1 = 23'b10011101110011010111110;
12'b001111001101: finv1 = 23'b10011101101110001001011;
12'b001111001110: finv1 = 23'b10011101101000111011001;
12'b001111001111: finv1 = 23'b10011101100011101101001;
12'b001111010000: finv1 = 23'b10011101011110011111001;
12'b001111010001: finv1 = 23'b10011101011001010001010;
12'b001111010010: finv1 = 23'b10011101010100000011100;
12'b001111010011: finv1 = 23'b10011101001110110110000;
12'b001111010100: finv1 = 23'b10011101001001101000100;
12'b001111010101: finv1 = 23'b10011101000100011011001;
12'b001111010110: finv1 = 23'b10011100111111001110000;
12'b001111010111: finv1 = 23'b10011100111010000000111;
12'b001111011000: finv1 = 23'b10011100110100110100000;
12'b001111011001: finv1 = 23'b10011100101111100111010;
12'b001111011010: finv1 = 23'b10011100101010011010100;
12'b001111011011: finv1 = 23'b10011100100101001110000;
12'b001111011100: finv1 = 23'b10011100100000000001101;
12'b001111011101: finv1 = 23'b10011100011010110101011;
12'b001111011110: finv1 = 23'b10011100010101101001010;
12'b001111011111: finv1 = 23'b10011100010000011101010;
12'b001111100000: finv1 = 23'b10011100001011010001010;
12'b001111100001: finv1 = 23'b10011100000110000101100;
12'b001111100010: finv1 = 23'b10011100000000111010000;
12'b001111100011: finv1 = 23'b10011011111011101110100;
12'b001111100100: finv1 = 23'b10011011110110100011001;
12'b001111100101: finv1 = 23'b10011011110001010111111;
12'b001111100110: finv1 = 23'b10011011101100001100110;
12'b001111100111: finv1 = 23'b10011011100111000001110;
12'b001111101000: finv1 = 23'b10011011100001110111000;
12'b001111101001: finv1 = 23'b10011011011100101100010;
12'b001111101010: finv1 = 23'b10011011010111100001101;
12'b001111101011: finv1 = 23'b10011011010010010111010;
12'b001111101100: finv1 = 23'b10011011001101001100111;
12'b001111101101: finv1 = 23'b10011011001000000010110;
12'b001111101110: finv1 = 23'b10011011000010111000101;
12'b001111101111: finv1 = 23'b10011010111101101110110;
12'b001111110000: finv1 = 23'b10011010111000100100111;
12'b001111110001: finv1 = 23'b10011010110011011011010;
12'b001111110010: finv1 = 23'b10011010101110010001110;
12'b001111110011: finv1 = 23'b10011010101001001000010;
12'b001111110100: finv1 = 23'b10011010100011111111000;
12'b001111110101: finv1 = 23'b10011010011110110101111;
12'b001111110110: finv1 = 23'b10011010011001101100111;
12'b001111110111: finv1 = 23'b10011010010100100011111;
12'b001111111000: finv1 = 23'b10011010001111011011001;
12'b001111111001: finv1 = 23'b10011010001010010010100;
12'b001111111010: finv1 = 23'b10011010000101001010000;
12'b001111111011: finv1 = 23'b10011010000000000001101;
12'b001111111100: finv1 = 23'b10011001111010111001011;
12'b001111111101: finv1 = 23'b10011001110101110001010;
12'b001111111110: finv1 = 23'b10011001110000101001010;
12'b001111111111: finv1 = 23'b10011001101011100001011;
12'b010000000000: finv1 = 23'b10011001100110011001101;
12'b010000000001: finv1 = 23'b10011001100001010010000;
12'b010000000010: finv1 = 23'b10011001011100001010100;
12'b010000000011: finv1 = 23'b10011001010111000011001;
12'b010000000100: finv1 = 23'b10011001010001111011111;
12'b010000000101: finv1 = 23'b10011001001100110100110;
12'b010000000110: finv1 = 23'b10011001000111101101111;
12'b010000000111: finv1 = 23'b10011001000010100111000;
12'b010000001000: finv1 = 23'b10011000111101100000010;
12'b010000001001: finv1 = 23'b10011000111000011001101;
12'b010000001010: finv1 = 23'b10011000110011010011010;
12'b010000001011: finv1 = 23'b10011000101110001100111;
12'b010000001100: finv1 = 23'b10011000101001000110101;
12'b010000001101: finv1 = 23'b10011000100100000000100;
12'b010000001110: finv1 = 23'b10011000011110111010101;
12'b010000001111: finv1 = 23'b10011000011001110100110;
12'b010000010000: finv1 = 23'b10011000010100101111000;
12'b010000010001: finv1 = 23'b10011000001111101001100;
12'b010000010010: finv1 = 23'b10011000001010100100000;
12'b010000010011: finv1 = 23'b10011000000101011110110;
12'b010000010100: finv1 = 23'b10011000000000011001100;
12'b010000010101: finv1 = 23'b10010111111011010100011;
12'b010000010110: finv1 = 23'b10010111110110001111100;
12'b010000010111: finv1 = 23'b10010111110001001010101;
12'b010000011000: finv1 = 23'b10010111101100000110000;
12'b010000011001: finv1 = 23'b10010111100111000001011;
12'b010000011010: finv1 = 23'b10010111100001111101000;
12'b010000011011: finv1 = 23'b10010111011100111000101;
12'b010000011100: finv1 = 23'b10010111010111110100100;
12'b010000011101: finv1 = 23'b10010111010010110000011;
12'b010000011110: finv1 = 23'b10010111001101101100100;
12'b010000011111: finv1 = 23'b10010111001000101000101;
12'b010000100000: finv1 = 23'b10010111000011100101000;
12'b010000100001: finv1 = 23'b10010110111110100001011;
12'b010000100010: finv1 = 23'b10010110111001011110000;
12'b010000100011: finv1 = 23'b10010110110100011010101;
12'b010000100100: finv1 = 23'b10010110101111010111100;
12'b010000100101: finv1 = 23'b10010110101010010100011;
12'b010000100110: finv1 = 23'b10010110100101010001100;
12'b010000100111: finv1 = 23'b10010110100000001110110;
12'b010000101000: finv1 = 23'b10010110011011001100000;
12'b010000101001: finv1 = 23'b10010110010110001001100;
12'b010000101010: finv1 = 23'b10010110010001000111000;
12'b010000101011: finv1 = 23'b10010110001100000100110;
12'b010000101100: finv1 = 23'b10010110000111000010100;
12'b010000101101: finv1 = 23'b10010110000010000000100;
12'b010000101110: finv1 = 23'b10010101111100111110100;
12'b010000101111: finv1 = 23'b10010101110111111100110;
12'b010000110000: finv1 = 23'b10010101110010111011000;
12'b010000110001: finv1 = 23'b10010101101101111001100;
12'b010000110010: finv1 = 23'b10010101101000111000000;
12'b010000110011: finv1 = 23'b10010101100011110110110;
12'b010000110100: finv1 = 23'b10010101011110110101100;
12'b010000110101: finv1 = 23'b10010101011001110100100;
12'b010000110110: finv1 = 23'b10010101010100110011100;
12'b010000110111: finv1 = 23'b10010101001111110010110;
12'b010000111000: finv1 = 23'b10010101001010110010000;
12'b010000111001: finv1 = 23'b10010101000101110001100;
12'b010000111010: finv1 = 23'b10010101000000110001000;
12'b010000111011: finv1 = 23'b10010100111011110000110;
12'b010000111100: finv1 = 23'b10010100110110110000100;
12'b010000111101: finv1 = 23'b10010100110001110000100;
12'b010000111110: finv1 = 23'b10010100101100110000100;
12'b010000111111: finv1 = 23'b10010100100111110000110;
12'b010001000000: finv1 = 23'b10010100100010110001000;
12'b010001000001: finv1 = 23'b10010100011101110001011;
12'b010001000010: finv1 = 23'b10010100011000110010000;
12'b010001000011: finv1 = 23'b10010100010011110010101;
12'b010001000100: finv1 = 23'b10010100001110110011011;
12'b010001000101: finv1 = 23'b10010100001001110100011;
12'b010001000110: finv1 = 23'b10010100000100110101011;
12'b010001000111: finv1 = 23'b10010011111111110110100;
12'b010001001000: finv1 = 23'b10010011111010110111111;
12'b010001001001: finv1 = 23'b10010011110101111001010;
12'b010001001010: finv1 = 23'b10010011110000111010110;
12'b010001001011: finv1 = 23'b10010011101011111100011;
12'b010001001100: finv1 = 23'b10010011100110111110001;
12'b010001001101: finv1 = 23'b10010011100010000000001;
12'b010001001110: finv1 = 23'b10010011011101000010001;
12'b010001001111: finv1 = 23'b10010011011000000100010;
12'b010001010000: finv1 = 23'b10010011010011000110100;
12'b010001010001: finv1 = 23'b10010011001110001000111;
12'b010001010010: finv1 = 23'b10010011001001001011011;
12'b010001010011: finv1 = 23'b10010011000100001110000;
12'b010001010100: finv1 = 23'b10010010111111010000110;
12'b010001010101: finv1 = 23'b10010010111010010011101;
12'b010001010110: finv1 = 23'b10010010110101010110101;
12'b010001010111: finv1 = 23'b10010010110000011001110;
12'b010001011000: finv1 = 23'b10010010101011011101000;
12'b010001011001: finv1 = 23'b10010010100110100000011;
12'b010001011010: finv1 = 23'b10010010100001100011111;
12'b010001011011: finv1 = 23'b10010010011100100111100;
12'b010001011100: finv1 = 23'b10010010010111101011001;
12'b010001011101: finv1 = 23'b10010010010010101111000;
12'b010001011110: finv1 = 23'b10010010001101110011000;
12'b010001011111: finv1 = 23'b10010010001000110111001;
12'b010001100000: finv1 = 23'b10010010000011111011010;
12'b010001100001: finv1 = 23'b10010001111110111111101;
12'b010001100010: finv1 = 23'b10010001111010000100001;
12'b010001100011: finv1 = 23'b10010001110101001000101;
12'b010001100100: finv1 = 23'b10010001110000001101011;
12'b010001100101: finv1 = 23'b10010001101011010010001;
12'b010001100110: finv1 = 23'b10010001100110010111001;
12'b010001100111: finv1 = 23'b10010001100001011100001;
12'b010001101000: finv1 = 23'b10010001011100100001011;
12'b010001101001: finv1 = 23'b10010001010111100110101;
12'b010001101010: finv1 = 23'b10010001010010101100000;
12'b010001101011: finv1 = 23'b10010001001101110001101;
12'b010001101100: finv1 = 23'b10010001001000110111010;
12'b010001101101: finv1 = 23'b10010001000011111101000;
12'b010001101110: finv1 = 23'b10010000111111000010111;
12'b010001101111: finv1 = 23'b10010000111010001000111;
12'b010001110000: finv1 = 23'b10010000110101001111001;
12'b010001110001: finv1 = 23'b10010000110000010101011;
12'b010001110010: finv1 = 23'b10010000101011011011110;
12'b010001110011: finv1 = 23'b10010000100110100010010;
12'b010001110100: finv1 = 23'b10010000100001101000111;
12'b010001110101: finv1 = 23'b10010000011100101111101;
12'b010001110110: finv1 = 23'b10010000010111110110011;
12'b010001110111: finv1 = 23'b10010000010010111101011;
12'b010001111000: finv1 = 23'b10010000001110000100100;
12'b010001111001: finv1 = 23'b10010000001001001011110;
12'b010001111010: finv1 = 23'b10010000000100010011000;
12'b010001111011: finv1 = 23'b10001111111111011010100;
12'b010001111100: finv1 = 23'b10001111111010100010001;
12'b010001111101: finv1 = 23'b10001111110101101001110;
12'b010001111110: finv1 = 23'b10001111110000110001101;
12'b010001111111: finv1 = 23'b10001111101011111001100;
12'b010010000000: finv1 = 23'b10001111100111000001100;
12'b010010000001: finv1 = 23'b10001111100010001001110;
12'b010010000010: finv1 = 23'b10001111011101010010000;
12'b010010000011: finv1 = 23'b10001111011000011010011;
12'b010010000100: finv1 = 23'b10001111010011100011000;
12'b010010000101: finv1 = 23'b10001111001110101011101;
12'b010010000110: finv1 = 23'b10001111001001110100011;
12'b010010000111: finv1 = 23'b10001111000100111101010;
12'b010010001000: finv1 = 23'b10001111000000000110010;
12'b010010001001: finv1 = 23'b10001110111011001111011;
12'b010010001010: finv1 = 23'b10001110110110011000101;
12'b010010001011: finv1 = 23'b10001110110001100010000;
12'b010010001100: finv1 = 23'b10001110101100101011011;
12'b010010001101: finv1 = 23'b10001110100111110101000;
12'b010010001110: finv1 = 23'b10001110100010111110110;
12'b010010001111: finv1 = 23'b10001110011110001000100;
12'b010010010000: finv1 = 23'b10001110011001010010100;
12'b010010010001: finv1 = 23'b10001110010100011100100;
12'b010010010010: finv1 = 23'b10001110001111100110110;
12'b010010010011: finv1 = 23'b10001110001010110001000;
12'b010010010100: finv1 = 23'b10001110000101111011011;
12'b010010010101: finv1 = 23'b10001110000001000110000;
12'b010010010110: finv1 = 23'b10001101111100010000101;
12'b010010010111: finv1 = 23'b10001101110111011011011;
12'b010010011000: finv1 = 23'b10001101110010100110010;
12'b010010011001: finv1 = 23'b10001101101101110001010;
12'b010010011010: finv1 = 23'b10001101101000111100011;
12'b010010011011: finv1 = 23'b10001101100100000111101;
12'b010010011100: finv1 = 23'b10001101011111010011000;
12'b010010011101: finv1 = 23'b10001101011010011110100;
12'b010010011110: finv1 = 23'b10001101010101101010000;
12'b010010011111: finv1 = 23'b10001101010000110101110;
12'b010010100000: finv1 = 23'b10001101001100000001100;
12'b010010100001: finv1 = 23'b10001101000111001101100;
12'b010010100010: finv1 = 23'b10001101000010011001100;
12'b010010100011: finv1 = 23'b10001100111101100101110;
12'b010010100100: finv1 = 23'b10001100111000110010000;
12'b010010100101: finv1 = 23'b10001100110011111110011;
12'b010010100110: finv1 = 23'b10001100101111001010111;
12'b010010100111: finv1 = 23'b10001100101010010111100;
12'b010010101000: finv1 = 23'b10001100100101100100010;
12'b010010101001: finv1 = 23'b10001100100000110001001;
12'b010010101010: finv1 = 23'b10001100011011111110001;
12'b010010101011: finv1 = 23'b10001100010111001011010;
12'b010010101100: finv1 = 23'b10001100010010011000100;
12'b010010101101: finv1 = 23'b10001100001101100101110;
12'b010010101110: finv1 = 23'b10001100001000110011010;
12'b010010101111: finv1 = 23'b10001100000100000000111;
12'b010010110000: finv1 = 23'b10001011111111001110100;
12'b010010110001: finv1 = 23'b10001011111010011100010;
12'b010010110010: finv1 = 23'b10001011110101101010010;
12'b010010110011: finv1 = 23'b10001011110000111000010;
12'b010010110100: finv1 = 23'b10001011101100000110011;
12'b010010110101: finv1 = 23'b10001011100111010100101;
12'b010010110110: finv1 = 23'b10001011100010100011000;
12'b010010110111: finv1 = 23'b10001011011101110001100;
12'b010010111000: finv1 = 23'b10001011011001000000001;
12'b010010111001: finv1 = 23'b10001011010100001110111;
12'b010010111010: finv1 = 23'b10001011001111011101101;
12'b010010111011: finv1 = 23'b10001011001010101100101;
12'b010010111100: finv1 = 23'b10001011000101111011101;
12'b010010111101: finv1 = 23'b10001011000001001010111;
12'b010010111110: finv1 = 23'b10001010111100011010001;
12'b010010111111: finv1 = 23'b10001010110111101001100;
12'b010011000000: finv1 = 23'b10001010110010111001000;
12'b010011000001: finv1 = 23'b10001010101110001000110;
12'b010011000010: finv1 = 23'b10001010101001011000100;
12'b010011000011: finv1 = 23'b10001010100100101000011;
12'b010011000100: finv1 = 23'b10001010011111111000010;
12'b010011000101: finv1 = 23'b10001010011011001000011;
12'b010011000110: finv1 = 23'b10001010010110011000101;
12'b010011000111: finv1 = 23'b10001010010001101000111;
12'b010011001000: finv1 = 23'b10001010001100111001011;
12'b010011001001: finv1 = 23'b10001010001000001001111;
12'b010011001010: finv1 = 23'b10001010000011011010101;
12'b010011001011: finv1 = 23'b10001001111110101011011;
12'b010011001100: finv1 = 23'b10001001111001111100010;
12'b010011001101: finv1 = 23'b10001001110101001101010;
12'b010011001110: finv1 = 23'b10001001110000011110011;
12'b010011001111: finv1 = 23'b10001001101011101111101;
12'b010011010000: finv1 = 23'b10001001100111000001000;
12'b010011010001: finv1 = 23'b10001001100010010010011;
12'b010011010010: finv1 = 23'b10001001011101100100000;
12'b010011010011: finv1 = 23'b10001001011000110101101;
12'b010011010100: finv1 = 23'b10001001010100000111100;
12'b010011010101: finv1 = 23'b10001001001111011001011;
12'b010011010110: finv1 = 23'b10001001001010101011011;
12'b010011010111: finv1 = 23'b10001001000101111101101;
12'b010011011000: finv1 = 23'b10001001000001001111111;
12'b010011011001: finv1 = 23'b10001000111100100010010;
12'b010011011010: finv1 = 23'b10001000110111110100101;
12'b010011011011: finv1 = 23'b10001000110011000111010;
12'b010011011100: finv1 = 23'b10001000101110011010000;
12'b010011011101: finv1 = 23'b10001000101001101100110;
12'b010011011110: finv1 = 23'b10001000100100111111110;
12'b010011011111: finv1 = 23'b10001000100000010010110;
12'b010011100000: finv1 = 23'b10001000011011100110000;
12'b010011100001: finv1 = 23'b10001000010110111001010;
12'b010011100010: finv1 = 23'b10001000010010001100101;
12'b010011100011: finv1 = 23'b10001000001101100000001;
12'b010011100100: finv1 = 23'b10001000001000110011110;
12'b010011100101: finv1 = 23'b10001000000100000111011;
12'b010011100110: finv1 = 23'b10000111111111011011010;
12'b010011100111: finv1 = 23'b10000111111010101111010;
12'b010011101000: finv1 = 23'b10000111110110000011010;
12'b010011101001: finv1 = 23'b10000111110001010111011;
12'b010011101010: finv1 = 23'b10000111101100101011110;
12'b010011101011: finv1 = 23'b10000111101000000000001;
12'b010011101100: finv1 = 23'b10000111100011010100101;
12'b010011101101: finv1 = 23'b10000111011110101001010;
12'b010011101110: finv1 = 23'b10000111011001111110000;
12'b010011101111: finv1 = 23'b10000111010101010010110;
12'b010011110000: finv1 = 23'b10000111010000100111110;
12'b010011110001: finv1 = 23'b10000111001011111100110;
12'b010011110010: finv1 = 23'b10000111000111010010000;
12'b010011110011: finv1 = 23'b10000111000010100111010;
12'b010011110100: finv1 = 23'b10000110111101111100101;
12'b010011110101: finv1 = 23'b10000110111001010010001;
12'b010011110110: finv1 = 23'b10000110110100100111110;
12'b010011110111: finv1 = 23'b10000110101111111101100;
12'b010011111000: finv1 = 23'b10000110101011010011011;
12'b010011111001: finv1 = 23'b10000110100110101001011;
12'b010011111010: finv1 = 23'b10000110100001111111011;
12'b010011111011: finv1 = 23'b10000110011101010101100;
12'b010011111100: finv1 = 23'b10000110011000101011111;
12'b010011111101: finv1 = 23'b10000110010100000010010;
12'b010011111110: finv1 = 23'b10000110001111011000110;
12'b010011111111: finv1 = 23'b10000110001010101111011;
12'b010100000000: finv1 = 23'b10000110000110000110001;
12'b010100000001: finv1 = 23'b10000110000001011100111;
12'b010100000010: finv1 = 23'b10000101111100110011111;
12'b010100000011: finv1 = 23'b10000101111000001011000;
12'b010100000100: finv1 = 23'b10000101110011100010001;
12'b010100000101: finv1 = 23'b10000101101110111001011;
12'b010100000110: finv1 = 23'b10000101101010010000110;
12'b010100000111: finv1 = 23'b10000101100101101000010;
12'b010100001000: finv1 = 23'b10000101100000111111111;
12'b010100001001: finv1 = 23'b10000101011100010111101;
12'b010100001010: finv1 = 23'b10000101010111101111100;
12'b010100001011: finv1 = 23'b10000101010011000111011;
12'b010100001100: finv1 = 23'b10000101001110011111100;
12'b010100001101: finv1 = 23'b10000101001001110111101;
12'b010100001110: finv1 = 23'b10000101000101001111111;
12'b010100001111: finv1 = 23'b10000101000000101000010;
12'b010100010000: finv1 = 23'b10000100111100000000110;
12'b010100010001: finv1 = 23'b10000100110111011001011;
12'b010100010010: finv1 = 23'b10000100110010110010001;
12'b010100010011: finv1 = 23'b10000100101110001010111;
12'b010100010100: finv1 = 23'b10000100101001100011111;
12'b010100010101: finv1 = 23'b10000100100100111100111;
12'b010100010110: finv1 = 23'b10000100100000010110000;
12'b010100010111: finv1 = 23'b10000100011011101111010;
12'b010100011000: finv1 = 23'b10000100010111001000101;
12'b010100011001: finv1 = 23'b10000100010010100010001;
12'b010100011010: finv1 = 23'b10000100001101111011110;
12'b010100011011: finv1 = 23'b10000100001001010101011;
12'b010100011100: finv1 = 23'b10000100000100101111001;
12'b010100011101: finv1 = 23'b10000100000000001001001;
12'b010100011110: finv1 = 23'b10000011111011100011001;
12'b010100011111: finv1 = 23'b10000011110110111101010;
12'b010100100000: finv1 = 23'b10000011110010010111100;
12'b010100100001: finv1 = 23'b10000011101101110001111;
12'b010100100010: finv1 = 23'b10000011101001001100010;
12'b010100100011: finv1 = 23'b10000011100100100110111;
12'b010100100100: finv1 = 23'b10000011100000000001100;
12'b010100100101: finv1 = 23'b10000011011011011100010;
12'b010100100110: finv1 = 23'b10000011010110110111001;
12'b010100100111: finv1 = 23'b10000011010010010010001;
12'b010100101000: finv1 = 23'b10000011001101101101010;
12'b010100101001: finv1 = 23'b10000011001001001000100;
12'b010100101010: finv1 = 23'b10000011000100100011111;
12'b010100101011: finv1 = 23'b10000010111111111111010;
12'b010100101100: finv1 = 23'b10000010111011011010110;
12'b010100101101: finv1 = 23'b10000010110110110110011;
12'b010100101110: finv1 = 23'b10000010110010010010001;
12'b010100101111: finv1 = 23'b10000010101101101110000;
12'b010100110000: finv1 = 23'b10000010101001001010000;
12'b010100110001: finv1 = 23'b10000010100100100110001;
12'b010100110010: finv1 = 23'b10000010100000000010010;
12'b010100110011: finv1 = 23'b10000010011011011110100;
12'b010100110100: finv1 = 23'b10000010010110111011000;
12'b010100110101: finv1 = 23'b10000010010010010111100;
12'b010100110110: finv1 = 23'b10000010001101110100001;
12'b010100110111: finv1 = 23'b10000010001001010000110;
12'b010100111000: finv1 = 23'b10000010000100101101101;
12'b010100111001: finv1 = 23'b10000010000000001010100;
12'b010100111010: finv1 = 23'b10000001111011100111101;
12'b010100111011: finv1 = 23'b10000001110111000100110;
12'b010100111100: finv1 = 23'b10000001110010100010000;
12'b010100111101: finv1 = 23'b10000001101101111111011;
12'b010100111110: finv1 = 23'b10000001101001011100111;
12'b010100111111: finv1 = 23'b10000001100100111010011;
12'b010101000000: finv1 = 23'b10000001100000011000001;
12'b010101000001: finv1 = 23'b10000001011011110101111;
12'b010101000010: finv1 = 23'b10000001010111010011110;
12'b010101000011: finv1 = 23'b10000001010010110001110;
12'b010101000100: finv1 = 23'b10000001001110001111111;
12'b010101000101: finv1 = 23'b10000001001001101110001;
12'b010101000110: finv1 = 23'b10000001000101001100011;
12'b010101000111: finv1 = 23'b10000001000000101010111;
12'b010101001000: finv1 = 23'b10000000111100001001011;
12'b010101001001: finv1 = 23'b10000000110111101000000;
12'b010101001010: finv1 = 23'b10000000110011000110110;
12'b010101001011: finv1 = 23'b10000000101110100101101;
12'b010101001100: finv1 = 23'b10000000101010000100101;
12'b010101001101: finv1 = 23'b10000000100101100011101;
12'b010101001110: finv1 = 23'b10000000100001000010111;
12'b010101001111: finv1 = 23'b10000000011100100010001;
12'b010101010000: finv1 = 23'b10000000011000000001100;
12'b010101010001: finv1 = 23'b10000000010011100001000;
12'b010101010010: finv1 = 23'b10000000001111000000101;
12'b010101010011: finv1 = 23'b10000000001010100000010;
12'b010101010100: finv1 = 23'b10000000000110000000001;
12'b010101010101: finv1 = 23'b10000000000001100000000;
12'b010101010110: finv1 = 23'b01111111111101000000000;
12'b010101010111: finv1 = 23'b01111111111000100000001;
12'b010101011000: finv1 = 23'b01111111110100000000011;
12'b010101011001: finv1 = 23'b01111111101111100000110;
12'b010101011010: finv1 = 23'b01111111101011000001001;
12'b010101011011: finv1 = 23'b01111111100110100001110;
12'b010101011100: finv1 = 23'b01111111100010000010011;
12'b010101011101: finv1 = 23'b01111111011101100011001;
12'b010101011110: finv1 = 23'b01111111011001000100000;
12'b010101011111: finv1 = 23'b01111111010100100100111;
12'b010101100000: finv1 = 23'b01111111010000000110000;
12'b010101100001: finv1 = 23'b01111111001011100111001;
12'b010101100010: finv1 = 23'b01111111000111001000100;
12'b010101100011: finv1 = 23'b01111111000010101001111;
12'b010101100100: finv1 = 23'b01111110111110001011011;
12'b010101100101: finv1 = 23'b01111110111001101100111;
12'b010101100110: finv1 = 23'b01111110110101001110101;
12'b010101100111: finv1 = 23'b01111110110000110000011;
12'b010101101000: finv1 = 23'b01111110101100010010010;
12'b010101101001: finv1 = 23'b01111110100111110100011;
12'b010101101010: finv1 = 23'b01111110100011010110100;
12'b010101101011: finv1 = 23'b01111110011110111000101;
12'b010101101100: finv1 = 23'b01111110011010011011000;
12'b010101101101: finv1 = 23'b01111110010101111101011;
12'b010101101110: finv1 = 23'b01111110010001100000000;
12'b010101101111: finv1 = 23'b01111110001101000010101;
12'b010101110000: finv1 = 23'b01111110001000100101011;
12'b010101110001: finv1 = 23'b01111110000100001000001;
12'b010101110010: finv1 = 23'b01111101111111101011001;
12'b010101110011: finv1 = 23'b01111101111011001110001;
12'b010101110100: finv1 = 23'b01111101110110110001011;
12'b010101110101: finv1 = 23'b01111101110010010100101;
12'b010101110110: finv1 = 23'b01111101101101111000000;
12'b010101110111: finv1 = 23'b01111101101001011011011;
12'b010101111000: finv1 = 23'b01111101100100111111000;
12'b010101111001: finv1 = 23'b01111101100000100010101;
12'b010101111010: finv1 = 23'b01111101011100000110011;
12'b010101111011: finv1 = 23'b01111101010111101010010;
12'b010101111100: finv1 = 23'b01111101010011001110010;
12'b010101111101: finv1 = 23'b01111101001110110010011;
12'b010101111110: finv1 = 23'b01111101001010010110101;
12'b010101111111: finv1 = 23'b01111101000101111010111;
12'b010110000000: finv1 = 23'b01111101000001011111010;
12'b010110000001: finv1 = 23'b01111100111101000011110;
12'b010110000010: finv1 = 23'b01111100111000101000011;
12'b010110000011: finv1 = 23'b01111100110100001101001;
12'b010110000100: finv1 = 23'b01111100101111110001111;
12'b010110000101: finv1 = 23'b01111100101011010110110;
12'b010110000110: finv1 = 23'b01111100100110111011110;
12'b010110000111: finv1 = 23'b01111100100010100000111;
12'b010110001000: finv1 = 23'b01111100011110000110001;
12'b010110001001: finv1 = 23'b01111100011001101011100;
12'b010110001010: finv1 = 23'b01111100010101010000111;
12'b010110001011: finv1 = 23'b01111100010000110110011;
12'b010110001100: finv1 = 23'b01111100001100011100000;
12'b010110001101: finv1 = 23'b01111100001000000001110;
12'b010110001110: finv1 = 23'b01111100000011100111101;
12'b010110001111: finv1 = 23'b01111011111111001101100;
12'b010110010000: finv1 = 23'b01111011111010110011101;
12'b010110010001: finv1 = 23'b01111011110110011001110;
12'b010110010010: finv1 = 23'b01111011110010000000000;
12'b010110010011: finv1 = 23'b01111011101101100110010;
12'b010110010100: finv1 = 23'b01111011101001001100110;
12'b010110010101: finv1 = 23'b01111011100100110011010;
12'b010110010110: finv1 = 23'b01111011100000011010000;
12'b010110010111: finv1 = 23'b01111011011100000000110;
12'b010110011000: finv1 = 23'b01111011010111100111100;
12'b010110011001: finv1 = 23'b01111011010011001110100;
12'b010110011010: finv1 = 23'b01111011001110110101100;
12'b010110011011: finv1 = 23'b01111011001010011100110;
12'b010110011100: finv1 = 23'b01111011000110000100000;
12'b010110011101: finv1 = 23'b01111011000001101011011;
12'b010110011110: finv1 = 23'b01111010111101010010110;
12'b010110011111: finv1 = 23'b01111010111000111010011;
12'b010110100000: finv1 = 23'b01111010110100100010000;
12'b010110100001: finv1 = 23'b01111010110000001001110;
12'b010110100010: finv1 = 23'b01111010101011110001101;
12'b010110100011: finv1 = 23'b01111010100111011001101;
12'b010110100100: finv1 = 23'b01111010100011000001110;
12'b010110100101: finv1 = 23'b01111010011110101001111;
12'b010110100110: finv1 = 23'b01111010011010010010001;
12'b010110100111: finv1 = 23'b01111010010101111010100;
12'b010110101000: finv1 = 23'b01111010010001100011000;
12'b010110101001: finv1 = 23'b01111010001101001011101;
12'b010110101010: finv1 = 23'b01111010001000110100010;
12'b010110101011: finv1 = 23'b01111010000100011101000;
12'b010110101100: finv1 = 23'b01111010000000000101111;
12'b010110101101: finv1 = 23'b01111001111011101110111;
12'b010110101110: finv1 = 23'b01111001110111011000000;
12'b010110101111: finv1 = 23'b01111001110011000001001;
12'b010110110000: finv1 = 23'b01111001101110101010011;
12'b010110110001: finv1 = 23'b01111001101010010011110;
12'b010110110010: finv1 = 23'b01111001100101111101010;
12'b010110110011: finv1 = 23'b01111001100001100110111;
12'b010110110100: finv1 = 23'b01111001011101010000100;
12'b010110110101: finv1 = 23'b01111001011000111010011;
12'b010110110110: finv1 = 23'b01111001010100100100010;
12'b010110110111: finv1 = 23'b01111001010000001110001;
12'b010110111000: finv1 = 23'b01111001001011111000010;
12'b010110111001: finv1 = 23'b01111001000111100010100;
12'b010110111010: finv1 = 23'b01111001000011001100110;
12'b010110111011: finv1 = 23'b01111000111110110111001;
12'b010110111100: finv1 = 23'b01111000111010100001101;
12'b010110111101: finv1 = 23'b01111000110110001100001;
12'b010110111110: finv1 = 23'b01111000110001110110111;
12'b010110111111: finv1 = 23'b01111000101101100001101;
12'b010111000000: finv1 = 23'b01111000101001001100100;
12'b010111000001: finv1 = 23'b01111000100100110111100;
12'b010111000010: finv1 = 23'b01111000100000100010100;
12'b010111000011: finv1 = 23'b01111000011100001101110;
12'b010111000100: finv1 = 23'b01111000010111111001000;
12'b010111000101: finv1 = 23'b01111000010011100100011;
12'b010111000110: finv1 = 23'b01111000001111001111111;
12'b010111000111: finv1 = 23'b01111000001010111011100;
12'b010111001000: finv1 = 23'b01111000000110100111001;
12'b010111001001: finv1 = 23'b01111000000010010010111;
12'b010111001010: finv1 = 23'b01110111111101111110110;
12'b010111001011: finv1 = 23'b01110111111001101010110;
12'b010111001100: finv1 = 23'b01110111110101010110110;
12'b010111001101: finv1 = 23'b01110111110001000011000;
12'b010111001110: finv1 = 23'b01110111101100101111010;
12'b010111001111: finv1 = 23'b01110111101000011011101;
12'b010111010000: finv1 = 23'b01110111100100001000001;
12'b010111010001: finv1 = 23'b01110111011111110100101;
12'b010111010010: finv1 = 23'b01110111011011100001010;
12'b010111010011: finv1 = 23'b01110111010111001110000;
12'b010111010100: finv1 = 23'b01110111010010111010111;
12'b010111010101: finv1 = 23'b01110111001110100111111;
12'b010111010110: finv1 = 23'b01110111001010010100111;
12'b010111010111: finv1 = 23'b01110111000110000010001;
12'b010111011000: finv1 = 23'b01110111000001101111011;
12'b010111011001: finv1 = 23'b01110110111101011100101;
12'b010111011010: finv1 = 23'b01110110111001001010001;
12'b010111011011: finv1 = 23'b01110110110100110111101;
12'b010111011100: finv1 = 23'b01110110110000100101011;
12'b010111011101: finv1 = 23'b01110110101100010011001;
12'b010111011110: finv1 = 23'b01110110101000000000111;
12'b010111011111: finv1 = 23'b01110110100011101110111;
12'b010111100000: finv1 = 23'b01110110011111011100111;
12'b010111100001: finv1 = 23'b01110110011011001011000;
12'b010111100010: finv1 = 23'b01110110010110111001010;
12'b010111100011: finv1 = 23'b01110110010010100111101;
12'b010111100100: finv1 = 23'b01110110001110010110000;
12'b010111100101: finv1 = 23'b01110110001010000100100;
12'b010111100110: finv1 = 23'b01110110000101110011001;
12'b010111100111: finv1 = 23'b01110110000001100001111;
12'b010111101000: finv1 = 23'b01110101111101010000110;
12'b010111101001: finv1 = 23'b01110101111000111111101;
12'b010111101010: finv1 = 23'b01110101110100101110101;
12'b010111101011: finv1 = 23'b01110101110000011101110;
12'b010111101100: finv1 = 23'b01110101101100001101000;
12'b010111101101: finv1 = 23'b01110101100111111100010;
12'b010111101110: finv1 = 23'b01110101100011101011101;
12'b010111101111: finv1 = 23'b01110101011111011011001;
12'b010111110000: finv1 = 23'b01110101011011001010110;
12'b010111110001: finv1 = 23'b01110101010110111010100;
12'b010111110010: finv1 = 23'b01110101010010101010010;
12'b010111110011: finv1 = 23'b01110101001110011010001;
12'b010111110100: finv1 = 23'b01110101001010001010001;
12'b010111110101: finv1 = 23'b01110101000101111010010;
12'b010111110110: finv1 = 23'b01110101000001101010011;
12'b010111110111: finv1 = 23'b01110100111101011010101;
12'b010111111000: finv1 = 23'b01110100111001001011000;
12'b010111111001: finv1 = 23'b01110100110100111011100;
12'b010111111010: finv1 = 23'b01110100110000101100000;
12'b010111111011: finv1 = 23'b01110100101100011100110;
12'b010111111100: finv1 = 23'b01110100101000001101100;
12'b010111111101: finv1 = 23'b01110100100011111110011;
12'b010111111110: finv1 = 23'b01110100011111101111010;
12'b010111111111: finv1 = 23'b01110100011011100000011;
12'b011000000000: finv1 = 23'b01110100010111010001100;
12'b011000000001: finv1 = 23'b01110100010011000010110;
12'b011000000010: finv1 = 23'b01110100001110110100000;
12'b011000000011: finv1 = 23'b01110100001010100101100;
12'b011000000100: finv1 = 23'b01110100000110010111000;
12'b011000000101: finv1 = 23'b01110100000010001000101;
12'b011000000110: finv1 = 23'b01110011111101111010011;
12'b011000000111: finv1 = 23'b01110011111001101100001;
12'b011000001000: finv1 = 23'b01110011110101011110000;
12'b011000001001: finv1 = 23'b01110011110001010000000;
12'b011000001010: finv1 = 23'b01110011101101000010001;
12'b011000001011: finv1 = 23'b01110011101000110100011;
12'b011000001100: finv1 = 23'b01110011100100100110101;
12'b011000001101: finv1 = 23'b01110011100000011001000;
12'b011000001110: finv1 = 23'b01110011011100001011100;
12'b011000001111: finv1 = 23'b01110011010111111110001;
12'b011000010000: finv1 = 23'b01110011010011110000110;
12'b011000010001: finv1 = 23'b01110011001111100011100;
12'b011000010010: finv1 = 23'b01110011001011010110011;
12'b011000010011: finv1 = 23'b01110011000111001001011;
12'b011000010100: finv1 = 23'b01110011000010111100011;
12'b011000010101: finv1 = 23'b01110010111110101111101;
12'b011000010110: finv1 = 23'b01110010111010100010111;
12'b011000010111: finv1 = 23'b01110010110110010110001;
12'b011000011000: finv1 = 23'b01110010110010001001101;
12'b011000011001: finv1 = 23'b01110010101101111101001;
12'b011000011010: finv1 = 23'b01110010101001110000110;
12'b011000011011: finv1 = 23'b01110010100101100100100;
12'b011000011100: finv1 = 23'b01110010100001011000010;
12'b011000011101: finv1 = 23'b01110010011101001100010;
12'b011000011110: finv1 = 23'b01110010011001000000010;
12'b011000011111: finv1 = 23'b01110010010100110100010;
12'b011000100000: finv1 = 23'b01110010010000101000100;
12'b011000100001: finv1 = 23'b01110010001100011100110;
12'b011000100010: finv1 = 23'b01110010001000010001001;
12'b011000100011: finv1 = 23'b01110010000100000101101;
12'b011000100100: finv1 = 23'b01110001111111111010010;
12'b011000100101: finv1 = 23'b01110001111011101110111;
12'b011000100110: finv1 = 23'b01110001110111100011101;
12'b011000100111: finv1 = 23'b01110001110011011000100;
12'b011000101000: finv1 = 23'b01110001101111001101100;
12'b011000101001: finv1 = 23'b01110001101011000010100;
12'b011000101010: finv1 = 23'b01110001100110110111101;
12'b011000101011: finv1 = 23'b01110001100010101100111;
12'b011000101100: finv1 = 23'b01110001011110100010001;
12'b011000101101: finv1 = 23'b01110001011010010111101;
12'b011000101110: finv1 = 23'b01110001010110001101001;
12'b011000101111: finv1 = 23'b01110001010010000010110;
12'b011000110000: finv1 = 23'b01110001001101111000011;
12'b011000110001: finv1 = 23'b01110001001001101110010;
12'b011000110010: finv1 = 23'b01110001000101100100001;
12'b011000110011: finv1 = 23'b01110001000001011010001;
12'b011000110100: finv1 = 23'b01110000111101010000001;
12'b011000110101: finv1 = 23'b01110000111001000110011;
12'b011000110110: finv1 = 23'b01110000110100111100101;
12'b011000110111: finv1 = 23'b01110000110000110011000;
12'b011000111000: finv1 = 23'b01110000101100101001011;
12'b011000111001: finv1 = 23'b01110000101000100000000;
12'b011000111010: finv1 = 23'b01110000100100010110101;
12'b011000111011: finv1 = 23'b01110000100000001101011;
12'b011000111100: finv1 = 23'b01110000011100000100001;
12'b011000111101: finv1 = 23'b01110000010111111011000;
12'b011000111110: finv1 = 23'b01110000010011110010001;
12'b011000111111: finv1 = 23'b01110000001111101001001;
12'b011001000000: finv1 = 23'b01110000001011100000011;
12'b011001000001: finv1 = 23'b01110000000111010111101;
12'b011001000010: finv1 = 23'b01110000000011001111000;
12'b011001000011: finv1 = 23'b01101111111111000110100;
12'b011001000100: finv1 = 23'b01101111111010111110001;
12'b011001000101: finv1 = 23'b01101111110110110101110;
12'b011001000110: finv1 = 23'b01101111110010101101100;
12'b011001000111: finv1 = 23'b01101111101110100101011;
12'b011001001000: finv1 = 23'b01101111101010011101010;
12'b011001001001: finv1 = 23'b01101111100110010101010;
12'b011001001010: finv1 = 23'b01101111100010001101011;
12'b011001001011: finv1 = 23'b01101111011110000101101;
12'b011001001100: finv1 = 23'b01101111011001111101111;
12'b011001001101: finv1 = 23'b01101111010101110110011;
12'b011001001110: finv1 = 23'b01101111010001101110111;
12'b011001001111: finv1 = 23'b01101111001101100111011;
12'b011001010000: finv1 = 23'b01101111001001100000001;
12'b011001010001: finv1 = 23'b01101111000101011000111;
12'b011001010010: finv1 = 23'b01101111000001010001110;
12'b011001010011: finv1 = 23'b01101110111101001010101;
12'b011001010100: finv1 = 23'b01101110111001000011110;
12'b011001010101: finv1 = 23'b01101110110100111100111;
12'b011001010110: finv1 = 23'b01101110110000110110001;
12'b011001010111: finv1 = 23'b01101110101100101111011;
12'b011001011000: finv1 = 23'b01101110101000101000111;
12'b011001011001: finv1 = 23'b01101110100100100010011;
12'b011001011010: finv1 = 23'b01101110100000011011111;
12'b011001011011: finv1 = 23'b01101110011100010101101;
12'b011001011100: finv1 = 23'b01101110011000001111011;
12'b011001011101: finv1 = 23'b01101110010100001001010;
12'b011001011110: finv1 = 23'b01101110010000000011010;
12'b011001011111: finv1 = 23'b01101110001011111101010;
12'b011001100000: finv1 = 23'b01101110000111110111011;
12'b011001100001: finv1 = 23'b01101110000011110001101;
12'b011001100010: finv1 = 23'b01101101111111101100000;
12'b011001100011: finv1 = 23'b01101101111011100110011;
12'b011001100100: finv1 = 23'b01101101110111100000111;
12'b011001100101: finv1 = 23'b01101101110011011011100;
12'b011001100110: finv1 = 23'b01101101101111010110010;
12'b011001100111: finv1 = 23'b01101101101011010001000;
12'b011001101000: finv1 = 23'b01101101100111001011111;
12'b011001101001: finv1 = 23'b01101101100011000110111;
12'b011001101010: finv1 = 23'b01101101011111000001111;
12'b011001101011: finv1 = 23'b01101101011010111101000;
12'b011001101100: finv1 = 23'b01101101010110111000010;
12'b011001101101: finv1 = 23'b01101101010010110011101;
12'b011001101110: finv1 = 23'b01101101001110101111000;
12'b011001101111: finv1 = 23'b01101101001010101010100;
12'b011001110000: finv1 = 23'b01101101000110100110001;
12'b011001110001: finv1 = 23'b01101101000010100001111;
12'b011001110010: finv1 = 23'b01101100111110011101101;
12'b011001110011: finv1 = 23'b01101100111010011001100;
12'b011001110100: finv1 = 23'b01101100110110010101100;
12'b011001110101: finv1 = 23'b01101100110010010001100;
12'b011001110110: finv1 = 23'b01101100101110001101101;
12'b011001110111: finv1 = 23'b01101100101010001001111;
12'b011001111000: finv1 = 23'b01101100100110000110010;
12'b011001111001: finv1 = 23'b01101100100010000010101;
12'b011001111010: finv1 = 23'b01101100011101111111001;
12'b011001111011: finv1 = 23'b01101100011001111011110;
12'b011001111100: finv1 = 23'b01101100010101111000100;
12'b011001111101: finv1 = 23'b01101100010001110101010;
12'b011001111110: finv1 = 23'b01101100001101110010001;
12'b011001111111: finv1 = 23'b01101100001001101111000;
12'b011010000000: finv1 = 23'b01101100000101101100001;
12'b011010000001: finv1 = 23'b01101100000001101001010;
12'b011010000010: finv1 = 23'b01101011111101100110100;
12'b011010000011: finv1 = 23'b01101011111001100011110;
12'b011010000100: finv1 = 23'b01101011110101100001001;
12'b011010000101: finv1 = 23'b01101011110001011110101;
12'b011010000110: finv1 = 23'b01101011101101011100010;
12'b011010000111: finv1 = 23'b01101011101001011001111;
12'b011010001000: finv1 = 23'b01101011100101010111110;
12'b011010001001: finv1 = 23'b01101011100001010101100;
12'b011010001010: finv1 = 23'b01101011011101010011100;
12'b011010001011: finv1 = 23'b01101011011001010001100;
12'b011010001100: finv1 = 23'b01101011010101001111101;
12'b011010001101: finv1 = 23'b01101011010001001101111;
12'b011010001110: finv1 = 23'b01101011001101001100001;
12'b011010001111: finv1 = 23'b01101011001001001010100;
12'b011010010000: finv1 = 23'b01101011000101001001000;
12'b011010010001: finv1 = 23'b01101011000001000111101;
12'b011010010010: finv1 = 23'b01101010111101000110010;
12'b011010010011: finv1 = 23'b01101010111001000101000;
12'b011010010100: finv1 = 23'b01101010110101000011111;
12'b011010010101: finv1 = 23'b01101010110001000010110;
12'b011010010110: finv1 = 23'b01101010101101000001110;
12'b011010010111: finv1 = 23'b01101010101001000000111;
12'b011010011000: finv1 = 23'b01101010100101000000001;
12'b011010011001: finv1 = 23'b01101010100000111111011;
12'b011010011010: finv1 = 23'b01101010011100111110110;
12'b011010011011: finv1 = 23'b01101010011000111110010;
12'b011010011100: finv1 = 23'b01101010010100111101110;
12'b011010011101: finv1 = 23'b01101010010000111101011;
12'b011010011110: finv1 = 23'b01101010001100111101001;
12'b011010011111: finv1 = 23'b01101010001000111100111;
12'b011010100000: finv1 = 23'b01101010000100111100111;
12'b011010100001: finv1 = 23'b01101010000000111100110;
12'b011010100010: finv1 = 23'b01101001111100111100111;
12'b011010100011: finv1 = 23'b01101001111000111101000;
12'b011010100100: finv1 = 23'b01101001110100111101010;
12'b011010100101: finv1 = 23'b01101001110000111101101;
12'b011010100110: finv1 = 23'b01101001101100111110001;
12'b011010100111: finv1 = 23'b01101001101000111110101;
12'b011010101000: finv1 = 23'b01101001100100111111010;
12'b011010101001: finv1 = 23'b01101001100000111111111;
12'b011010101010: finv1 = 23'b01101001011101000000101;
12'b011010101011: finv1 = 23'b01101001011001000001100;
12'b011010101100: finv1 = 23'b01101001010101000010100;
12'b011010101101: finv1 = 23'b01101001010001000011100;
12'b011010101110: finv1 = 23'b01101001001101000100110;
12'b011010101111: finv1 = 23'b01101001001001000101111;
12'b011010110000: finv1 = 23'b01101001000101000111010;
12'b011010110001: finv1 = 23'b01101001000001001000101;
12'b011010110010: finv1 = 23'b01101000111101001010001;
12'b011010110011: finv1 = 23'b01101000111001001011101;
12'b011010110100: finv1 = 23'b01101000110101001101011;
12'b011010110101: finv1 = 23'b01101000110001001111001;
12'b011010110110: finv1 = 23'b01101000101101010000111;
12'b011010110111: finv1 = 23'b01101000101001010010111;
12'b011010111000: finv1 = 23'b01101000100101010100111;
12'b011010111001: finv1 = 23'b01101000100001010111000;
12'b011010111010: finv1 = 23'b01101000011101011001001;
12'b011010111011: finv1 = 23'b01101000011001011011011;
12'b011010111100: finv1 = 23'b01101000010101011101110;
12'b011010111101: finv1 = 23'b01101000010001100000010;
12'b011010111110: finv1 = 23'b01101000001101100010110;
12'b011010111111: finv1 = 23'b01101000001001100101011;
12'b011011000000: finv1 = 23'b01101000000101101000001;
12'b011011000001: finv1 = 23'b01101000000001101010111;
12'b011011000010: finv1 = 23'b01100111111101101101110;
12'b011011000011: finv1 = 23'b01100111111001110000110;
12'b011011000100: finv1 = 23'b01100111110101110011110;
12'b011011000101: finv1 = 23'b01100111110001110110111;
12'b011011000110: finv1 = 23'b01100111101101111010001;
12'b011011000111: finv1 = 23'b01100111101001111101100;
12'b011011001000: finv1 = 23'b01100111100110000000111;
12'b011011001001: finv1 = 23'b01100111100010000100011;
12'b011011001010: finv1 = 23'b01100111011110001000000;
12'b011011001011: finv1 = 23'b01100111011010001011101;
12'b011011001100: finv1 = 23'b01100111010110001111011;
12'b011011001101: finv1 = 23'b01100111010010010011010;
12'b011011001110: finv1 = 23'b01100111001110010111001;
12'b011011001111: finv1 = 23'b01100111001010011011001;
12'b011011010000: finv1 = 23'b01100111000110011111010;
12'b011011010001: finv1 = 23'b01100111000010100011011;
12'b011011010010: finv1 = 23'b01100110111110100111101;
12'b011011010011: finv1 = 23'b01100110111010101100000;
12'b011011010100: finv1 = 23'b01100110110110110000100;
12'b011011010101: finv1 = 23'b01100110110010110101000;
12'b011011010110: finv1 = 23'b01100110101110111001101;
12'b011011010111: finv1 = 23'b01100110101010111110010;
12'b011011011000: finv1 = 23'b01100110100111000011001;
12'b011011011001: finv1 = 23'b01100110100011000111111;
12'b011011011010: finv1 = 23'b01100110011111001100111;
12'b011011011011: finv1 = 23'b01100110011011010001111;
12'b011011011100: finv1 = 23'b01100110010111010111000;
12'b011011011101: finv1 = 23'b01100110010011011100010;
12'b011011011110: finv1 = 23'b01100110001111100001101;
12'b011011011111: finv1 = 23'b01100110001011100111000;
12'b011011100000: finv1 = 23'b01100110000111101100011;
12'b011011100001: finv1 = 23'b01100110000011110010000;
12'b011011100010: finv1 = 23'b01100101111111110111101;
12'b011011100011: finv1 = 23'b01100101111011111101011;
12'b011011100100: finv1 = 23'b01100101111000000011001;
12'b011011100101: finv1 = 23'b01100101110100001001000;
12'b011011100110: finv1 = 23'b01100101110000001111000;
12'b011011100111: finv1 = 23'b01100101101100010101001;
12'b011011101000: finv1 = 23'b01100101101000011011010;
12'b011011101001: finv1 = 23'b01100101100100100001100;
12'b011011101010: finv1 = 23'b01100101100000100111110;
12'b011011101011: finv1 = 23'b01100101011100101110010;
12'b011011101100: finv1 = 23'b01100101011000110100110;
12'b011011101101: finv1 = 23'b01100101010100111011010;
12'b011011101110: finv1 = 23'b01100101010001000010000;
12'b011011101111: finv1 = 23'b01100101001101001000110;
12'b011011110000: finv1 = 23'b01100101001001001111100;
12'b011011110001: finv1 = 23'b01100101000101010110100;
12'b011011110010: finv1 = 23'b01100101000001011101100;
12'b011011110011: finv1 = 23'b01100100111101100100100;
12'b011011110100: finv1 = 23'b01100100111001101011110;
12'b011011110101: finv1 = 23'b01100100110101110011000;
12'b011011110110: finv1 = 23'b01100100110001111010010;
12'b011011110111: finv1 = 23'b01100100101110000001110;
12'b011011111000: finv1 = 23'b01100100101010001001010;
12'b011011111001: finv1 = 23'b01100100100110010000111;
12'b011011111010: finv1 = 23'b01100100100010011000100;
12'b011011111011: finv1 = 23'b01100100011110100000010;
12'b011011111100: finv1 = 23'b01100100011010101000001;
12'b011011111101: finv1 = 23'b01100100010110110000000;
12'b011011111110: finv1 = 23'b01100100010010111000001;
12'b011011111111: finv1 = 23'b01100100001111000000001;
12'b011100000000: finv1 = 23'b01100100001011001000011;
12'b011100000001: finv1 = 23'b01100100000111010000101;
12'b011100000010: finv1 = 23'b01100100000011011001000;
12'b011100000011: finv1 = 23'b01100011111111100001011;
12'b011100000100: finv1 = 23'b01100011111011101001111;
12'b011100000101: finv1 = 23'b01100011110111110010100;
12'b011100000110: finv1 = 23'b01100011110011111011010;
12'b011100000111: finv1 = 23'b01100011110000000100000;
12'b011100001000: finv1 = 23'b01100011101100001100111;
12'b011100001001: finv1 = 23'b01100011101000010101110;
12'b011100001010: finv1 = 23'b01100011100100011110111;
12'b011100001011: finv1 = 23'b01100011100000100111111;
12'b011100001100: finv1 = 23'b01100011011100110001001;
12'b011100001101: finv1 = 23'b01100011011000111010011;
12'b011100001110: finv1 = 23'b01100011010101000011110;
12'b011100001111: finv1 = 23'b01100011010001001101010;
12'b011100010000: finv1 = 23'b01100011001101010110110;
12'b011100010001: finv1 = 23'b01100011001001100000011;
12'b011100010010: finv1 = 23'b01100011000101101010000;
12'b011100010011: finv1 = 23'b01100011000001110011110;
12'b011100010100: finv1 = 23'b01100010111101111101101;
12'b011100010101: finv1 = 23'b01100010111010000111101;
12'b011100010110: finv1 = 23'b01100010110110010001101;
12'b011100010111: finv1 = 23'b01100010110010011011110;
12'b011100011000: finv1 = 23'b01100010101110100101111;
12'b011100011001: finv1 = 23'b01100010101010110000010;
12'b011100011010: finv1 = 23'b01100010100110111010101;
12'b011100011011: finv1 = 23'b01100010100011000101000;
12'b011100011100: finv1 = 23'b01100010011111001111100;
12'b011100011101: finv1 = 23'b01100010011011011010001;
12'b011100011110: finv1 = 23'b01100010010111100100111;
12'b011100011111: finv1 = 23'b01100010010011101111101;
12'b011100100000: finv1 = 23'b01100010001111111010100;
12'b011100100001: finv1 = 23'b01100010001100000101011;
12'b011100100010: finv1 = 23'b01100010001000010000011;
12'b011100100011: finv1 = 23'b01100010000100011011100;
12'b011100100100: finv1 = 23'b01100010000000100110110;
12'b011100100101: finv1 = 23'b01100001111100110010000;
12'b011100100110: finv1 = 23'b01100001111000111101011;
12'b011100100111: finv1 = 23'b01100001110101001000110;
12'b011100101000: finv1 = 23'b01100001110001010100010;
12'b011100101001: finv1 = 23'b01100001101101011111111;
12'b011100101010: finv1 = 23'b01100001101001101011101;
12'b011100101011: finv1 = 23'b01100001100101110111011;
12'b011100101100: finv1 = 23'b01100001100010000011010;
12'b011100101101: finv1 = 23'b01100001011110001111001;
12'b011100101110: finv1 = 23'b01100001011010011011001;
12'b011100101111: finv1 = 23'b01100001010110100111010;
12'b011100110000: finv1 = 23'b01100001010010110011011;
12'b011100110001: finv1 = 23'b01100001001110111111101;
12'b011100110010: finv1 = 23'b01100001001011001100000;
12'b011100110011: finv1 = 23'b01100001000111011000011;
12'b011100110100: finv1 = 23'b01100001000011100100111;
12'b011100110101: finv1 = 23'b01100000111111110001100;
12'b011100110110: finv1 = 23'b01100000111011111110010;
12'b011100110111: finv1 = 23'b01100000111000001011000;
12'b011100111000: finv1 = 23'b01100000110100010111110;
12'b011100111001: finv1 = 23'b01100000110000100100110;
12'b011100111010: finv1 = 23'b01100000101100110001101;
12'b011100111011: finv1 = 23'b01100000101000111110110;
12'b011100111100: finv1 = 23'b01100000100101001011111;
12'b011100111101: finv1 = 23'b01100000100001011001001;
12'b011100111110: finv1 = 23'b01100000011101100110100;
12'b011100111111: finv1 = 23'b01100000011001110011111;
12'b011101000000: finv1 = 23'b01100000010110000001011;
12'b011101000001: finv1 = 23'b01100000010010001111000;
12'b011101000010: finv1 = 23'b01100000001110011100101;
12'b011101000011: finv1 = 23'b01100000001010101010011;
12'b011101000100: finv1 = 23'b01100000000110111000001;
12'b011101000101: finv1 = 23'b01100000000011000110000;
12'b011101000110: finv1 = 23'b01011111111111010100000;
12'b011101000111: finv1 = 23'b01011111111011100010000;
12'b011101001000: finv1 = 23'b01011111110111110000010;
12'b011101001001: finv1 = 23'b01011111110011111110011;
12'b011101001010: finv1 = 23'b01011111110000001100110;
12'b011101001011: finv1 = 23'b01011111101100011011001;
12'b011101001100: finv1 = 23'b01011111101000101001100;
12'b011101001101: finv1 = 23'b01011111100100111000001;
12'b011101001110: finv1 = 23'b01011111100001000110110;
12'b011101001111: finv1 = 23'b01011111011101010101011;
12'b011101010000: finv1 = 23'b01011111011001100100010;
12'b011101010001: finv1 = 23'b01011111010101110011001;
12'b011101010010: finv1 = 23'b01011111010010000010000;
12'b011101010011: finv1 = 23'b01011111001110010001000;
12'b011101010100: finv1 = 23'b01011111001010100000001;
12'b011101010101: finv1 = 23'b01011111000110101111011;
12'b011101010110: finv1 = 23'b01011111000010111110101;
12'b011101010111: finv1 = 23'b01011110111111001110000;
12'b011101011000: finv1 = 23'b01011110111011011101011;
12'b011101011001: finv1 = 23'b01011110110111101100111;
12'b011101011010: finv1 = 23'b01011110110011111100100;
12'b011101011011: finv1 = 23'b01011110110000001100001;
12'b011101011100: finv1 = 23'b01011110101100011011111;
12'b011101011101: finv1 = 23'b01011110101000101011110;
12'b011101011110: finv1 = 23'b01011110100100111011101;
12'b011101011111: finv1 = 23'b01011110100001001011101;
12'b011101100000: finv1 = 23'b01011110011101011011110;
12'b011101100001: finv1 = 23'b01011110011001101011111;
12'b011101100010: finv1 = 23'b01011110010101111100001;
12'b011101100011: finv1 = 23'b01011110010010001100011;
12'b011101100100: finv1 = 23'b01011110001110011100111;
12'b011101100101: finv1 = 23'b01011110001010101101010;
12'b011101100110: finv1 = 23'b01011110000110111101111;
12'b011101100111: finv1 = 23'b01011110000011001110100;
12'b011101101000: finv1 = 23'b01011101111111011111010;
12'b011101101001: finv1 = 23'b01011101111011110000000;
12'b011101101010: finv1 = 23'b01011101111000000000111;
12'b011101101011: finv1 = 23'b01011101110100010001110;
12'b011101101100: finv1 = 23'b01011101110000100010111;
12'b011101101101: finv1 = 23'b01011101101100110100000;
12'b011101101110: finv1 = 23'b01011101101001000101001;
12'b011101101111: finv1 = 23'b01011101100101010110011;
12'b011101110000: finv1 = 23'b01011101100001100111110;
12'b011101110001: finv1 = 23'b01011101011101111001010;
12'b011101110010: finv1 = 23'b01011101011010001010110;
12'b011101110011: finv1 = 23'b01011101010110011100010;
12'b011101110100: finv1 = 23'b01011101010010101110000;
12'b011101110101: finv1 = 23'b01011101001110111111110;
12'b011101110110: finv1 = 23'b01011101001011010001100;
12'b011101110111: finv1 = 23'b01011101000111100011100;
12'b011101111000: finv1 = 23'b01011101000011110101011;
12'b011101111001: finv1 = 23'b01011101000000000111100;
12'b011101111010: finv1 = 23'b01011100111100011001101;
12'b011101111011: finv1 = 23'b01011100111000101011111;
12'b011101111100: finv1 = 23'b01011100110100111110001;
12'b011101111101: finv1 = 23'b01011100110001010000100;
12'b011101111110: finv1 = 23'b01011100101101100011000;
12'b011101111111: finv1 = 23'b01011100101001110101100;
12'b011110000000: finv1 = 23'b01011100100110001000001;
12'b011110000001: finv1 = 23'b01011100100010011010111;
12'b011110000010: finv1 = 23'b01011100011110101101101;
12'b011110000011: finv1 = 23'b01011100011011000000100;
12'b011110000100: finv1 = 23'b01011100010111010011011;
12'b011110000101: finv1 = 23'b01011100010011100110100;
12'b011110000110: finv1 = 23'b01011100001111111001100;
12'b011110000111: finv1 = 23'b01011100001100001100110;
12'b011110001000: finv1 = 23'b01011100001000100000000;
12'b011110001001: finv1 = 23'b01011100000100110011010;
12'b011110001010: finv1 = 23'b01011100000001000110110;
12'b011110001011: finv1 = 23'b01011011111101011010001;
12'b011110001100: finv1 = 23'b01011011111001101101110;
12'b011110001101: finv1 = 23'b01011011110110000001011;
12'b011110001110: finv1 = 23'b01011011110010010101001;
12'b011110001111: finv1 = 23'b01011011101110101000111;
12'b011110010000: finv1 = 23'b01011011101010111100110;
12'b011110010001: finv1 = 23'b01011011100111010000110;
12'b011110010010: finv1 = 23'b01011011100011100100110;
12'b011110010011: finv1 = 23'b01011011011111111000111;
12'b011110010100: finv1 = 23'b01011011011100001101001;
12'b011110010101: finv1 = 23'b01011011011000100001011;
12'b011110010110: finv1 = 23'b01011011010100110101101;
12'b011110010111: finv1 = 23'b01011011010001001010001;
12'b011110011000: finv1 = 23'b01011011001101011110101;
12'b011110011001: finv1 = 23'b01011011001001110011001;
12'b011110011010: finv1 = 23'b01011011000110000111111;
12'b011110011011: finv1 = 23'b01011011000010011100101;
12'b011110011100: finv1 = 23'b01011010111110110001011;
12'b011110011101: finv1 = 23'b01011010111011000110010;
12'b011110011110: finv1 = 23'b01011010110111011011010;
12'b011110011111: finv1 = 23'b01011010110011110000010;
12'b011110100000: finv1 = 23'b01011010110000000101011;
12'b011110100001: finv1 = 23'b01011010101100011010101;
12'b011110100010: finv1 = 23'b01011010101000101111111;
12'b011110100011: finv1 = 23'b01011010100101000101010;
12'b011110100100: finv1 = 23'b01011010100001011010110;
12'b011110100101: finv1 = 23'b01011010011101110000010;
12'b011110100110: finv1 = 23'b01011010011010000101110;
12'b011110100111: finv1 = 23'b01011010010110011011100;
12'b011110101000: finv1 = 23'b01011010010010110001010;
12'b011110101001: finv1 = 23'b01011010001111000111000;
12'b011110101010: finv1 = 23'b01011010001011011100111;
12'b011110101011: finv1 = 23'b01011010000111110010111;
12'b011110101100: finv1 = 23'b01011010000100001001000;
12'b011110101101: finv1 = 23'b01011010000000011111001;
12'b011110101110: finv1 = 23'b01011001111100110101010;
12'b011110101111: finv1 = 23'b01011001111001001011101;
12'b011110110000: finv1 = 23'b01011001110101100010000;
12'b011110110001: finv1 = 23'b01011001110001111000011;
12'b011110110010: finv1 = 23'b01011001101110001110111;
12'b011110110011: finv1 = 23'b01011001101010100101100;
12'b011110110100: finv1 = 23'b01011001100110111100001;
12'b011110110101: finv1 = 23'b01011001100011010010111;
12'b011110110110: finv1 = 23'b01011001011111101001110;
12'b011110110111: finv1 = 23'b01011001011100000000101;
12'b011110111000: finv1 = 23'b01011001011000010111101;
12'b011110111001: finv1 = 23'b01011001010100101110101;
12'b011110111010: finv1 = 23'b01011001010001000101110;
12'b011110111011: finv1 = 23'b01011001001101011101000;
12'b011110111100: finv1 = 23'b01011001001001110100010;
12'b011110111101: finv1 = 23'b01011001000110001011101;
12'b011110111110: finv1 = 23'b01011001000010100011001;
12'b011110111111: finv1 = 23'b01011000111110111010101;
12'b011111000000: finv1 = 23'b01011000111011010010010;
12'b011111000001: finv1 = 23'b01011000110111101001111;
12'b011111000010: finv1 = 23'b01011000110100000001101;
12'b011111000011: finv1 = 23'b01011000110000011001011;
12'b011111000100: finv1 = 23'b01011000101100110001011;
12'b011111000101: finv1 = 23'b01011000101001001001010;
12'b011111000110: finv1 = 23'b01011000100101100001011;
12'b011111000111: finv1 = 23'b01011000100001111001100;
12'b011111001000: finv1 = 23'b01011000011110010001101;
12'b011111001001: finv1 = 23'b01011000011010101010000;
12'b011111001010: finv1 = 23'b01011000010111000010010;
12'b011111001011: finv1 = 23'b01011000010011011010110;
12'b011111001100: finv1 = 23'b01011000001111110011010;
12'b011111001101: finv1 = 23'b01011000001100001011110;
12'b011111001110: finv1 = 23'b01011000001000100100100;
12'b011111001111: finv1 = 23'b01011000000100111101010;
12'b011111010000: finv1 = 23'b01011000000001010110000;
12'b011111010001: finv1 = 23'b01010111111101101110111;
12'b011111010010: finv1 = 23'b01010111111010000111111;
12'b011111010011: finv1 = 23'b01010111110110100000111;
12'b011111010100: finv1 = 23'b01010111110010111010000;
12'b011111010101: finv1 = 23'b01010111101111010011001;
12'b011111010110: finv1 = 23'b01010111101011101100100;
12'b011111010111: finv1 = 23'b01010111101000000101110;
12'b011111011000: finv1 = 23'b01010111100100011111010;
12'b011111011001: finv1 = 23'b01010111100000111000110;
12'b011111011010: finv1 = 23'b01010111011101010010010;
12'b011111011011: finv1 = 23'b01010111011001101011111;
12'b011111011100: finv1 = 23'b01010111010110000101101;
12'b011111011101: finv1 = 23'b01010111010010011111011;
12'b011111011110: finv1 = 23'b01010111001110111001010;
12'b011111011111: finv1 = 23'b01010111001011010011010;
12'b011111100000: finv1 = 23'b01010111000111101101010;
12'b011111100001: finv1 = 23'b01010111000100000111011;
12'b011111100010: finv1 = 23'b01010111000000100001100;
12'b011111100011: finv1 = 23'b01010110111100111011110;
12'b011111100100: finv1 = 23'b01010110111001010110000;
12'b011111100101: finv1 = 23'b01010110110101110000100;
12'b011111100110: finv1 = 23'b01010110110010001010111;
12'b011111100111: finv1 = 23'b01010110101110100101100;
12'b011111101000: finv1 = 23'b01010110101011000000001;
12'b011111101001: finv1 = 23'b01010110100111011010110;
12'b011111101010: finv1 = 23'b01010110100011110101100;
12'b011111101011: finv1 = 23'b01010110100000010000011;
12'b011111101100: finv1 = 23'b01010110011100101011010;
12'b011111101101: finv1 = 23'b01010110011001000110010;
12'b011111101110: finv1 = 23'b01010110010101100001011;
12'b011111101111: finv1 = 23'b01010110010001111100100;
12'b011111110000: finv1 = 23'b01010110001110010111110;
12'b011111110001: finv1 = 23'b01010110001010110011000;
12'b011111110010: finv1 = 23'b01010110000111001110011;
12'b011111110011: finv1 = 23'b01010110000011101001111;
12'b011111110100: finv1 = 23'b01010110000000000101011;
12'b011111110101: finv1 = 23'b01010101111100100000111;
12'b011111110110: finv1 = 23'b01010101111000111100101;
12'b011111110111: finv1 = 23'b01010101110101011000011;
12'b011111111000: finv1 = 23'b01010101110001110100001;
12'b011111111001: finv1 = 23'b01010101101110010000000;
12'b011111111010: finv1 = 23'b01010101101010101100000;
12'b011111111011: finv1 = 23'b01010101100111001000000;
12'b011111111100: finv1 = 23'b01010101100011100100001;
12'b011111111101: finv1 = 23'b01010101100000000000011;
12'b011111111110: finv1 = 23'b01010101011100011100101;
12'b011111111111: finv1 = 23'b01010101011000111000111;
12'b100000000000: finv1 = 23'b01010101010101010101011;
12'b100000000001: finv1 = 23'b01010101010001110001111;
12'b100000000010: finv1 = 23'b01010101001110001110011;
12'b100000000011: finv1 = 23'b01010101001010101011000;
12'b100000000100: finv1 = 23'b01010101000111000111110;
12'b100000000101: finv1 = 23'b01010101000011100100100;
12'b100000000110: finv1 = 23'b01010101000000000001011;
12'b100000000111: finv1 = 23'b01010100111100011110010;
12'b100000001000: finv1 = 23'b01010100111000111011010;
12'b100000001001: finv1 = 23'b01010100110101011000011;
12'b100000001010: finv1 = 23'b01010100110001110101100;
12'b100000001011: finv1 = 23'b01010100101110010010110;
12'b100000001100: finv1 = 23'b01010100101010110000000;
12'b100000001101: finv1 = 23'b01010100100111001101011;
12'b100000001110: finv1 = 23'b01010100100011101010110;
12'b100000001111: finv1 = 23'b01010100100000001000011;
12'b100000010000: finv1 = 23'b01010100011100100101111;
12'b100000010001: finv1 = 23'b01010100011001000011101;
12'b100000010010: finv1 = 23'b01010100010101100001010;
12'b100000010011: finv1 = 23'b01010100010001111111001;
12'b100000010100: finv1 = 23'b01010100001110011101000;
12'b100000010101: finv1 = 23'b01010100001010111011000;
12'b100000010110: finv1 = 23'b01010100000111011001000;
12'b100000010111: finv1 = 23'b01010100000011110111001;
12'b100000011000: finv1 = 23'b01010100000000010101010;
12'b100000011001: finv1 = 23'b01010011111100110011100;
12'b100000011010: finv1 = 23'b01010011111001010001111;
12'b100000011011: finv1 = 23'b01010011110101110000010;
12'b100000011100: finv1 = 23'b01010011110010001110101;
12'b100000011101: finv1 = 23'b01010011101110101101010;
12'b100000011110: finv1 = 23'b01010011101011001011111;
12'b100000011111: finv1 = 23'b01010011100111101010100;
12'b100000100000: finv1 = 23'b01010011100100001001010;
12'b100000100001: finv1 = 23'b01010011100000101000001;
12'b100000100010: finv1 = 23'b01010011011101000111000;
12'b100000100011: finv1 = 23'b01010011011001100110000;
12'b100000100100: finv1 = 23'b01010011010110000101000;
12'b100000100101: finv1 = 23'b01010011010010100100001;
12'b100000100110: finv1 = 23'b01010011001111000011011;
12'b100000100111: finv1 = 23'b01010011001011100010101;
12'b100000101000: finv1 = 23'b01010011001000000010000;
12'b100000101001: finv1 = 23'b01010011000100100001011;
12'b100000101010: finv1 = 23'b01010011000001000000111;
12'b100000101011: finv1 = 23'b01010010111101100000100;
12'b100000101100: finv1 = 23'b01010010111010000000001;
12'b100000101101: finv1 = 23'b01010010110110011111110;
12'b100000101110: finv1 = 23'b01010010110010111111101;
12'b100000101111: finv1 = 23'b01010010101111011111011;
12'b100000110000: finv1 = 23'b01010010101011111111011;
12'b100000110001: finv1 = 23'b01010010101000011111011;
12'b100000110010: finv1 = 23'b01010010100100111111011;
12'b100000110011: finv1 = 23'b01010010100001011111100;
12'b100000110100: finv1 = 23'b01010010011101111111110;
12'b100000110101: finv1 = 23'b01010010011010100000000;
12'b100000110110: finv1 = 23'b01010010010111000000011;
12'b100000110111: finv1 = 23'b01010010010011100000111;
12'b100000111000: finv1 = 23'b01010010010000000001011;
12'b100000111001: finv1 = 23'b01010010001100100001111;
12'b100000111010: finv1 = 23'b01010010001001000010100;
12'b100000111011: finv1 = 23'b01010010000101100011010;
12'b100000111100: finv1 = 23'b01010010000010000100000;
12'b100000111101: finv1 = 23'b01010001111110100100111;
12'b100000111110: finv1 = 23'b01010001111011000101111;
12'b100000111111: finv1 = 23'b01010001110111100110111;
12'b100001000000: finv1 = 23'b01010001110100000111111;
12'b100001000001: finv1 = 23'b01010001110000101001001;
12'b100001000010: finv1 = 23'b01010001101101001010010;
12'b100001000011: finv1 = 23'b01010001101001101011101;
12'b100001000100: finv1 = 23'b01010001100110001101000;
12'b100001000101: finv1 = 23'b01010001100010101110011;
12'b100001000110: finv1 = 23'b01010001011111001111111;
12'b100001000111: finv1 = 23'b01010001011011110001100;
12'b100001001000: finv1 = 23'b01010001011000010011001;
12'b100001001001: finv1 = 23'b01010001010100110100111;
12'b100001001010: finv1 = 23'b01010001010001010110101;
12'b100001001011: finv1 = 23'b01010001001101111000100;
12'b100001001100: finv1 = 23'b01010001001010011010011;
12'b100001001101: finv1 = 23'b01010001000110111100011;
12'b100001001110: finv1 = 23'b01010001000011011110100;
12'b100001001111: finv1 = 23'b01010001000000000000101;
12'b100001010000: finv1 = 23'b01010000111100100010111;
12'b100001010001: finv1 = 23'b01010000111001000101001;
12'b100001010010: finv1 = 23'b01010000110101100111100;
12'b100001010011: finv1 = 23'b01010000110010001010000;
12'b100001010100: finv1 = 23'b01010000101110101100100;
12'b100001010101: finv1 = 23'b01010000101011001111000;
12'b100001010110: finv1 = 23'b01010000100111110001110;
12'b100001010111: finv1 = 23'b01010000100100010100011;
12'b100001011000: finv1 = 23'b01010000100000110111010;
12'b100001011001: finv1 = 23'b01010000011101011010001;
12'b100001011010: finv1 = 23'b01010000011001111101000;
12'b100001011011: finv1 = 23'b01010000010110100000000;
12'b100001011100: finv1 = 23'b01010000010011000011001;
12'b100001011101: finv1 = 23'b01010000001111100110010;
12'b100001011110: finv1 = 23'b01010000001100001001100;
12'b100001011111: finv1 = 23'b01010000001000101100110;
12'b100001100000: finv1 = 23'b01010000000101010000001;
12'b100001100001: finv1 = 23'b01010000000001110011100;
12'b100001100010: finv1 = 23'b01001111111110010111000;
12'b100001100011: finv1 = 23'b01001111111010111010101;
12'b100001100100: finv1 = 23'b01001111110111011110010;
12'b100001100101: finv1 = 23'b01001111110100000001111;
12'b100001100110: finv1 = 23'b01001111110000100101110;
12'b100001100111: finv1 = 23'b01001111101101001001100;
12'b100001101000: finv1 = 23'b01001111101001101101100;
12'b100001101001: finv1 = 23'b01001111100110010001100;
12'b100001101010: finv1 = 23'b01001111100010110101100;
12'b100001101011: finv1 = 23'b01001111011111011001101;
12'b100001101100: finv1 = 23'b01001111011011111101111;
12'b100001101101: finv1 = 23'b01001111011000100010001;
12'b100001101110: finv1 = 23'b01001111010101000110100;
12'b100001101111: finv1 = 23'b01001111010001101010111;
12'b100001110000: finv1 = 23'b01001111001110001111011;
12'b100001110001: finv1 = 23'b01001111001010110100000;
12'b100001110010: finv1 = 23'b01001111000111011000101;
12'b100001110011: finv1 = 23'b01001111000011111101010;
12'b100001110100: finv1 = 23'b01001111000000100010000;
12'b100001110101: finv1 = 23'b01001110111101000110111;
12'b100001110110: finv1 = 23'b01001110111001101011110;
12'b100001110111: finv1 = 23'b01001110110110010000110;
12'b100001111000: finv1 = 23'b01001110110010110101110;
12'b100001111001: finv1 = 23'b01001110101111011010111;
12'b100001111010: finv1 = 23'b01001110101100000000001;
12'b100001111011: finv1 = 23'b01001110101000100101011;
12'b100001111100: finv1 = 23'b01001110100101001010101;
12'b100001111101: finv1 = 23'b01001110100001110000000;
12'b100001111110: finv1 = 23'b01001110011110010101100;
12'b100001111111: finv1 = 23'b01001110011010111011000;
12'b100010000000: finv1 = 23'b01001110010111100000101;
12'b100010000001: finv1 = 23'b01001110010100000110011;
12'b100010000010: finv1 = 23'b01001110010000101100001;
12'b100010000011: finv1 = 23'b01001110001101010001111;
12'b100010000100: finv1 = 23'b01001110001001110111110;
12'b100010000101: finv1 = 23'b01001110000110011101110;
12'b100010000110: finv1 = 23'b01001110000011000011110;
12'b100010000111: finv1 = 23'b01001101111111101001111;
12'b100010001000: finv1 = 23'b01001101111100010000000;
12'b100010001001: finv1 = 23'b01001101111000110110010;
12'b100010001010: finv1 = 23'b01001101110101011100100;
12'b100010001011: finv1 = 23'b01001101110010000010111;
12'b100010001100: finv1 = 23'b01001101101110101001010;
12'b100010001101: finv1 = 23'b01001101101011001111111;
12'b100010001110: finv1 = 23'b01001101100111110110011;
12'b100010001111: finv1 = 23'b01001101100100011101000;
12'b100010010000: finv1 = 23'b01001101100001000011110;
12'b100010010001: finv1 = 23'b01001101011101101010100;
12'b100010010010: finv1 = 23'b01001101011010010001011;
12'b100010010011: finv1 = 23'b01001101010110111000010;
12'b100010010100: finv1 = 23'b01001101010011011111010;
12'b100010010101: finv1 = 23'b01001101010000000110011;
12'b100010010110: finv1 = 23'b01001101001100101101100;
12'b100010010111: finv1 = 23'b01001101001001010100101;
12'b100010011000: finv1 = 23'b01001101000101111011111;
12'b100010011001: finv1 = 23'b01001101000010100011010;
12'b100010011010: finv1 = 23'b01001100111111001010101;
12'b100010011011: finv1 = 23'b01001100111011110010001;
12'b100010011100: finv1 = 23'b01001100111000011001101;
12'b100010011101: finv1 = 23'b01001100110101000001010;
12'b100010011110: finv1 = 23'b01001100110001101001000;
12'b100010011111: finv1 = 23'b01001100101110010000110;
12'b100010100000: finv1 = 23'b01001100101010111000100;
12'b100010100001: finv1 = 23'b01001100100111100000011;
12'b100010100010: finv1 = 23'b01001100100100001000011;
12'b100010100011: finv1 = 23'b01001100100000110000011;
12'b100010100100: finv1 = 23'b01001100011101011000100;
12'b100010100101: finv1 = 23'b01001100011010000000101;
12'b100010100110: finv1 = 23'b01001100010110101000111;
12'b100010100111: finv1 = 23'b01001100010011010001001;
12'b100010101000: finv1 = 23'b01001100001111111001100;
12'b100010101001: finv1 = 23'b01001100001100100010000;
12'b100010101010: finv1 = 23'b01001100001001001010100;
12'b100010101011: finv1 = 23'b01001100000101110011000;
12'b100010101100: finv1 = 23'b01001100000010011011101;
12'b100010101101: finv1 = 23'b01001011111111000100011;
12'b100010101110: finv1 = 23'b01001011111011101101001;
12'b100010101111: finv1 = 23'b01001011111000010110000;
12'b100010110000: finv1 = 23'b01001011110100111110111;
12'b100010110001: finv1 = 23'b01001011110001100111111;
12'b100010110010: finv1 = 23'b01001011101110010000111;
12'b100010110011: finv1 = 23'b01001011101010111010000;
12'b100010110100: finv1 = 23'b01001011100111100011001;
12'b100010110101: finv1 = 23'b01001011100100001100011;
12'b100010110110: finv1 = 23'b01001011100000110101110;
12'b100010110111: finv1 = 23'b01001011011101011111001;
12'b100010111000: finv1 = 23'b01001011011010001000101;
12'b100010111001: finv1 = 23'b01001011010110110010001;
12'b100010111010: finv1 = 23'b01001011010011011011101;
12'b100010111011: finv1 = 23'b01001011010000000101011;
12'b100010111100: finv1 = 23'b01001011001100101111000;
12'b100010111101: finv1 = 23'b01001011001001011000111;
12'b100010111110: finv1 = 23'b01001011000110000010110;
12'b100010111111: finv1 = 23'b01001011000010101100101;
12'b100011000000: finv1 = 23'b01001010111111010110101;
12'b100011000001: finv1 = 23'b01001010111100000000101;
12'b100011000010: finv1 = 23'b01001010111000101010111;
12'b100011000011: finv1 = 23'b01001010110101010101000;
12'b100011000100: finv1 = 23'b01001010110001111111010;
12'b100011000101: finv1 = 23'b01001010101110101001101;
12'b100011000110: finv1 = 23'b01001010101011010100000;
12'b100011000111: finv1 = 23'b01001010100111111110100;
12'b100011001000: finv1 = 23'b01001010100100101001000;
12'b100011001001: finv1 = 23'b01001010100001010011101;
12'b100011001010: finv1 = 23'b01001010011101111110010;
12'b100011001011: finv1 = 23'b01001010011010101001000;
12'b100011001100: finv1 = 23'b01001010010111010011110;
12'b100011001101: finv1 = 23'b01001010010011111110101;
12'b100011001110: finv1 = 23'b01001010010000101001101;
12'b100011001111: finv1 = 23'b01001010001101010100101;
12'b100011010000: finv1 = 23'b01001010001001111111101;
12'b100011010001: finv1 = 23'b01001010000110101010111;
12'b100011010010: finv1 = 23'b01001010000011010110000;
12'b100011010011: finv1 = 23'b01001010000000000001010;
12'b100011010100: finv1 = 23'b01001001111100101100101;
12'b100011010101: finv1 = 23'b01001001111001011000000;
12'b100011010110: finv1 = 23'b01001001110110000011100;
12'b100011010111: finv1 = 23'b01001001110010101111000;
12'b100011011000: finv1 = 23'b01001001101111011010101;
12'b100011011001: finv1 = 23'b01001001101100000110011;
12'b100011011010: finv1 = 23'b01001001101000110010000;
12'b100011011011: finv1 = 23'b01001001100101011101111;
12'b100011011100: finv1 = 23'b01001001100010001001110;
12'b100011011101: finv1 = 23'b01001001011110110101101;
12'b100011011110: finv1 = 23'b01001001011011100001101;
12'b100011011111: finv1 = 23'b01001001011000001101110;
12'b100011100000: finv1 = 23'b01001001010100111001111;
12'b100011100001: finv1 = 23'b01001001010001100110001;
12'b100011100010: finv1 = 23'b01001001001110010010011;
12'b100011100011: finv1 = 23'b01001001001010111110110;
12'b100011100100: finv1 = 23'b01001001000111101011001;
12'b100011100101: finv1 = 23'b01001001000100010111101;
12'b100011100110: finv1 = 23'b01001001000001000100001;
12'b100011100111: finv1 = 23'b01001000111101110000110;
12'b100011101000: finv1 = 23'b01001000111010011101011;
12'b100011101001: finv1 = 23'b01001000110111001010001;
12'b100011101010: finv1 = 23'b01001000110011110110111;
12'b100011101011: finv1 = 23'b01001000110000100011110;
12'b100011101100: finv1 = 23'b01001000101101010000110;
12'b100011101101: finv1 = 23'b01001000101001111101110;
12'b100011101110: finv1 = 23'b01001000100110101010110;
12'b100011101111: finv1 = 23'b01001000100011010111111;
12'b100011110000: finv1 = 23'b01001000100000000101001;
12'b100011110001: finv1 = 23'b01001000011100110010011;
12'b100011110010: finv1 = 23'b01001000011001011111110;
12'b100011110011: finv1 = 23'b01001000010110001101001;
12'b100011110100: finv1 = 23'b01001000010010111010101;
12'b100011110101: finv1 = 23'b01001000001111101000001;
12'b100011110110: finv1 = 23'b01001000001100010101110;
12'b100011110111: finv1 = 23'b01001000001001000011011;
12'b100011111000: finv1 = 23'b01001000000101110001001;
12'b100011111001: finv1 = 23'b01001000000010011110111;
12'b100011111010: finv1 = 23'b01000111111111001100110;
12'b100011111011: finv1 = 23'b01000111111011111010101;
12'b100011111100: finv1 = 23'b01000111111000101000101;
12'b100011111101: finv1 = 23'b01000111110101010110110;
12'b100011111110: finv1 = 23'b01000111110010000100111;
12'b100011111111: finv1 = 23'b01000111101110110011000;
12'b100100000000: finv1 = 23'b01000111101011100001010;
12'b100100000001: finv1 = 23'b01000111101000001111101;
12'b100100000010: finv1 = 23'b01000111100100111110000;
12'b100100000011: finv1 = 23'b01000111100001101100011;
12'b100100000100: finv1 = 23'b01000111011110011011000;
12'b100100000101: finv1 = 23'b01000111011011001001100;
12'b100100000110: finv1 = 23'b01000111010111111000001;
12'b100100000111: finv1 = 23'b01000111010100100110111;
12'b100100001000: finv1 = 23'b01000111010001010101101;
12'b100100001001: finv1 = 23'b01000111001110000100100;
12'b100100001010: finv1 = 23'b01000111001010110011011;
12'b100100001011: finv1 = 23'b01000111000111100010011;
12'b100100001100: finv1 = 23'b01000111000100010001011;
12'b100100001101: finv1 = 23'b01000111000001000000100;
12'b100100001110: finv1 = 23'b01000110111101101111101;
12'b100100001111: finv1 = 23'b01000110111010011110111;
12'b100100010000: finv1 = 23'b01000110110111001110010;
12'b100100010001: finv1 = 23'b01000110110011111101101;
12'b100100010010: finv1 = 23'b01000110110000101101000;
12'b100100010011: finv1 = 23'b01000110101101011100100;
12'b100100010100: finv1 = 23'b01000110101010001100000;
12'b100100010101: finv1 = 23'b01000110100110111011101;
12'b100100010110: finv1 = 23'b01000110100011101011011;
12'b100100010111: finv1 = 23'b01000110100000011011001;
12'b100100011000: finv1 = 23'b01000110011101001010111;
12'b100100011001: finv1 = 23'b01000110011001111010110;
12'b100100011010: finv1 = 23'b01000110010110101010110;
12'b100100011011: finv1 = 23'b01000110010011011010110;
12'b100100011100: finv1 = 23'b01000110010000001010111;
12'b100100011101: finv1 = 23'b01000110001100111011000;
12'b100100011110: finv1 = 23'b01000110001001101011001;
12'b100100011111: finv1 = 23'b01000110000110011011100;
12'b100100100000: finv1 = 23'b01000110000011001011110;
12'b100100100001: finv1 = 23'b01000101111111111100001;
12'b100100100010: finv1 = 23'b01000101111100101100101;
12'b100100100011: finv1 = 23'b01000101111001011101001;
12'b100100100100: finv1 = 23'b01000101110110001101110;
12'b100100100101: finv1 = 23'b01000101110010111110011;
12'b100100100110: finv1 = 23'b01000101101111101111001;
12'b100100100111: finv1 = 23'b01000101101100011111111;
12'b100100101000: finv1 = 23'b01000101101001010000110;
12'b100100101001: finv1 = 23'b01000101100110000001110;
12'b100100101010: finv1 = 23'b01000101100010110010101;
12'b100100101011: finv1 = 23'b01000101011111100011110;
12'b100100101100: finv1 = 23'b01000101011100010100111;
12'b100100101101: finv1 = 23'b01000101011001000110000;
12'b100100101110: finv1 = 23'b01000101010101110111010;
12'b100100101111: finv1 = 23'b01000101010010101000100;
12'b100100110000: finv1 = 23'b01000101001111011001111;
12'b100100110001: finv1 = 23'b01000101001100001011011;
12'b100100110010: finv1 = 23'b01000101001000111100110;
12'b100100110011: finv1 = 23'b01000101000101101110011;
12'b100100110100: finv1 = 23'b01000101000010100000000;
12'b100100110101: finv1 = 23'b01000100111111010001101;
12'b100100110110: finv1 = 23'b01000100111100000011011;
12'b100100110111: finv1 = 23'b01000100111000110101010;
12'b100100111000: finv1 = 23'b01000100110101100111001;
12'b100100111001: finv1 = 23'b01000100110010011001000;
12'b100100111010: finv1 = 23'b01000100101111001011000;
12'b100100111011: finv1 = 23'b01000100101011111101001;
12'b100100111100: finv1 = 23'b01000100101000101111010;
12'b100100111101: finv1 = 23'b01000100100101100001011;
12'b100100111110: finv1 = 23'b01000100100010010011110;
12'b100100111111: finv1 = 23'b01000100011111000110000;
12'b100101000000: finv1 = 23'b01000100011011111000011;
12'b100101000001: finv1 = 23'b01000100011000101010111;
12'b100101000010: finv1 = 23'b01000100010101011101011;
12'b100101000011: finv1 = 23'b01000100010010001111111;
12'b100101000100: finv1 = 23'b01000100001111000010101;
12'b100101000101: finv1 = 23'b01000100001011110101010;
12'b100101000110: finv1 = 23'b01000100001000101000000;
12'b100101000111: finv1 = 23'b01000100000101011010111;
12'b100101001000: finv1 = 23'b01000100000010001101110;
12'b100101001001: finv1 = 23'b01000011111111000000110;
12'b100101001010: finv1 = 23'b01000011111011110011110;
12'b100101001011: finv1 = 23'b01000011111000100110111;
12'b100101001100: finv1 = 23'b01000011110101011010000;
12'b100101001101: finv1 = 23'b01000011110010001101001;
12'b100101001110: finv1 = 23'b01000011101111000000100;
12'b100101001111: finv1 = 23'b01000011101011110011110;
12'b100101010000: finv1 = 23'b01000011101000100111010;
12'b100101010001: finv1 = 23'b01000011100101011010101;
12'b100101010010: finv1 = 23'b01000011100010001110001;
12'b100101010011: finv1 = 23'b01000011011111000001110;
12'b100101010100: finv1 = 23'b01000011011011110101011;
12'b100101010101: finv1 = 23'b01000011011000101001001;
12'b100101010110: finv1 = 23'b01000011010101011100111;
12'b100101010111: finv1 = 23'b01000011010010010000110;
12'b100101011000: finv1 = 23'b01000011001111000100101;
12'b100101011001: finv1 = 23'b01000011001011111000101;
12'b100101011010: finv1 = 23'b01000011001000101100101;
12'b100101011011: finv1 = 23'b01000011000101100000110;
12'b100101011100: finv1 = 23'b01000011000010010100111;
12'b100101011101: finv1 = 23'b01000010111111001001001;
12'b100101011110: finv1 = 23'b01000010111011111101011;
12'b100101011111: finv1 = 23'b01000010111000110001110;
12'b100101100000: finv1 = 23'b01000010110101100110001;
12'b100101100001: finv1 = 23'b01000010110010011010101;
12'b100101100010: finv1 = 23'b01000010101111001111001;
12'b100101100011: finv1 = 23'b01000010101100000011110;
12'b100101100100: finv1 = 23'b01000010101000111000011;
12'b100101100101: finv1 = 23'b01000010100101101101001;
12'b100101100110: finv1 = 23'b01000010100010100001111;
12'b100101100111: finv1 = 23'b01000010011111010110110;
12'b100101101000: finv1 = 23'b01000010011100001011101;
12'b100101101001: finv1 = 23'b01000010011001000000101;
12'b100101101010: finv1 = 23'b01000010010101110101101;
12'b100101101011: finv1 = 23'b01000010010010101010110;
12'b100101101100: finv1 = 23'b01000010001111011111111;
12'b100101101101: finv1 = 23'b01000010001100010101001;
12'b100101101110: finv1 = 23'b01000010001001001010011;
12'b100101101111: finv1 = 23'b01000010000101111111110;
12'b100101110000: finv1 = 23'b01000010000010110101001;
12'b100101110001: finv1 = 23'b01000001111111101010101;
12'b100101110010: finv1 = 23'b01000001111100100000001;
12'b100101110011: finv1 = 23'b01000001111001010101110;
12'b100101110100: finv1 = 23'b01000001110110001011011;
12'b100101110101: finv1 = 23'b01000001110011000001001;
12'b100101110110: finv1 = 23'b01000001101111110110111;
12'b100101110111: finv1 = 23'b01000001101100101100110;
12'b100101111000: finv1 = 23'b01000001101001100010101;
12'b100101111001: finv1 = 23'b01000001100110011000101;
12'b100101111010: finv1 = 23'b01000001100011001110101;
12'b100101111011: finv1 = 23'b01000001100000000100110;
12'b100101111100: finv1 = 23'b01000001011100111010111;
12'b100101111101: finv1 = 23'b01000001011001110001001;
12'b100101111110: finv1 = 23'b01000001010110100111011;
12'b100101111111: finv1 = 23'b01000001010011011101101;
12'b100110000000: finv1 = 23'b01000001010000010100001;
12'b100110000001: finv1 = 23'b01000001001101001010100;
12'b100110000010: finv1 = 23'b01000001001010000001000;
12'b100110000011: finv1 = 23'b01000001000110110111101;
12'b100110000100: finv1 = 23'b01000001000011101110010;
12'b100110000101: finv1 = 23'b01000001000000100101000;
12'b100110000110: finv1 = 23'b01000000111101011011110;
12'b100110000111: finv1 = 23'b01000000111010010010101;
12'b100110001000: finv1 = 23'b01000000110111001001100;
12'b100110001001: finv1 = 23'b01000000110100000000011;
12'b100110001010: finv1 = 23'b01000000110000110111100;
12'b100110001011: finv1 = 23'b01000000101101101110100;
12'b100110001100: finv1 = 23'b01000000101010100101101;
12'b100110001101: finv1 = 23'b01000000100111011100111;
12'b100110001110: finv1 = 23'b01000000100100010100001;
12'b100110001111: finv1 = 23'b01000000100001001011011;
12'b100110010000: finv1 = 23'b01000000011110000010111;
12'b100110010001: finv1 = 23'b01000000011010111010010;
12'b100110010010: finv1 = 23'b01000000010111110001110;
12'b100110010011: finv1 = 23'b01000000010100101001011;
12'b100110010100: finv1 = 23'b01000000010001100001000;
12'b100110010101: finv1 = 23'b01000000001110011000101;
12'b100110010110: finv1 = 23'b01000000001011010000011;
12'b100110010111: finv1 = 23'b01000000001000001000010;
12'b100110011000: finv1 = 23'b01000000000101000000001;
12'b100110011001: finv1 = 23'b01000000000001111000000;
12'b100110011010: finv1 = 23'b00111111111110110000000;
12'b100110011011: finv1 = 23'b00111111111011101000000;
12'b100110011100: finv1 = 23'b00111111111000100000001;
12'b100110011101: finv1 = 23'b00111111110101011000011;
12'b100110011110: finv1 = 23'b00111111110010010000101;
12'b100110011111: finv1 = 23'b00111111101111001000111;
12'b100110100000: finv1 = 23'b00111111101100000001010;
12'b100110100001: finv1 = 23'b00111111101000111001101;
12'b100110100010: finv1 = 23'b00111111100101110010001;
12'b100110100011: finv1 = 23'b00111111100010101010110;
12'b100110100100: finv1 = 23'b00111111011111100011010;
12'b100110100101: finv1 = 23'b00111111011100011100000;
12'b100110100110: finv1 = 23'b00111111011001010100101;
12'b100110100111: finv1 = 23'b00111111010110001101100;
12'b100110101000: finv1 = 23'b00111111010011000110011;
12'b100110101001: finv1 = 23'b00111111001111111111010;
12'b100110101010: finv1 = 23'b00111111001100111000010;
12'b100110101011: finv1 = 23'b00111111001001110001010;
12'b100110101100: finv1 = 23'b00111111000110101010010;
12'b100110101101: finv1 = 23'b00111111000011100011100;
12'b100110101110: finv1 = 23'b00111111000000011100101;
12'b100110101111: finv1 = 23'b00111110111101010101111;
12'b100110110000: finv1 = 23'b00111110111010001111010;
12'b100110110001: finv1 = 23'b00111110110111001000101;
12'b100110110010: finv1 = 23'b00111110110100000010001;
12'b100110110011: finv1 = 23'b00111110110000111011101;
12'b100110110100: finv1 = 23'b00111110101101110101001;
12'b100110110101: finv1 = 23'b00111110101010101110111;
12'b100110110110: finv1 = 23'b00111110100111101000100;
12'b100110110111: finv1 = 23'b00111110100100100010010;
12'b100110111000: finv1 = 23'b00111110100001011100001;
12'b100110111001: finv1 = 23'b00111110011110010110000;
12'b100110111010: finv1 = 23'b00111110011011001111111;
12'b100110111011: finv1 = 23'b00111110011000001001111;
12'b100110111100: finv1 = 23'b00111110010101000011111;
12'b100110111101: finv1 = 23'b00111110010001111110000;
12'b100110111110: finv1 = 23'b00111110001110111000010;
12'b100110111111: finv1 = 23'b00111110001011110010100;
12'b100111000000: finv1 = 23'b00111110001000101100110;
12'b100111000001: finv1 = 23'b00111110000101100111001;
12'b100111000010: finv1 = 23'b00111110000010100001100;
12'b100111000011: finv1 = 23'b00111101111111011100000;
12'b100111000100: finv1 = 23'b00111101111100010110100;
12'b100111000101: finv1 = 23'b00111101111001010001001;
12'b100111000110: finv1 = 23'b00111101110110001011110;
12'b100111000111: finv1 = 23'b00111101110011000110100;
12'b100111001000: finv1 = 23'b00111101110000000001010;
12'b100111001001: finv1 = 23'b00111101101100111100001;
12'b100111001010: finv1 = 23'b00111101101001110111000;
12'b100111001011: finv1 = 23'b00111101100110110001111;
12'b100111001100: finv1 = 23'b00111101100011101100111;
12'b100111001101: finv1 = 23'b00111101100000101000000;
12'b100111001110: finv1 = 23'b00111101011101100011001;
12'b100111001111: finv1 = 23'b00111101011010011110011;
12'b100111010000: finv1 = 23'b00111101010111011001101;
12'b100111010001: finv1 = 23'b00111101010100010100111;
12'b100111010010: finv1 = 23'b00111101010001010000010;
12'b100111010011: finv1 = 23'b00111101001110001011101;
12'b100111010100: finv1 = 23'b00111101001011000111001;
12'b100111010101: finv1 = 23'b00111101001000000010110;
12'b100111010110: finv1 = 23'b00111101000100111110011;
12'b100111010111: finv1 = 23'b00111101000001111010000;
12'b100111011000: finv1 = 23'b00111100111110110101110;
12'b100111011001: finv1 = 23'b00111100111011110001100;
12'b100111011010: finv1 = 23'b00111100111000101101011;
12'b100111011011: finv1 = 23'b00111100110101101001010;
12'b100111011100: finv1 = 23'b00111100110010100101010;
12'b100111011101: finv1 = 23'b00111100101111100001010;
12'b100111011110: finv1 = 23'b00111100101100011101010;
12'b100111011111: finv1 = 23'b00111100101001011001100;
12'b100111100000: finv1 = 23'b00111100100110010101101;
12'b100111100001: finv1 = 23'b00111100100011010001111;
12'b100111100010: finv1 = 23'b00111100100000001110010;
12'b100111100011: finv1 = 23'b00111100011101001010101;
12'b100111100100: finv1 = 23'b00111100011010000111000;
12'b100111100101: finv1 = 23'b00111100010111000011100;
12'b100111100110: finv1 = 23'b00111100010100000000001;
12'b100111100111: finv1 = 23'b00111100010000111100110;
12'b100111101000: finv1 = 23'b00111100001101111001011;
12'b100111101001: finv1 = 23'b00111100001010110110001;
12'b100111101010: finv1 = 23'b00111100000111110010111;
12'b100111101011: finv1 = 23'b00111100000100101111110;
12'b100111101100: finv1 = 23'b00111100000001101100101;
12'b100111101101: finv1 = 23'b00111011111110101001101;
12'b100111101110: finv1 = 23'b00111011111011100110101;
12'b100111101111: finv1 = 23'b00111011111000100011110;
12'b100111110000: finv1 = 23'b00111011110101100000111;
12'b100111110001: finv1 = 23'b00111011110010011110000;
12'b100111110010: finv1 = 23'b00111011101111011011010;
12'b100111110011: finv1 = 23'b00111011101100011000101;
12'b100111110100: finv1 = 23'b00111011101001010110000;
12'b100111110101: finv1 = 23'b00111011100110010011011;
12'b100111110110: finv1 = 23'b00111011100011010000111;
12'b100111110111: finv1 = 23'b00111011100000001110100;
12'b100111111000: finv1 = 23'b00111011011101001100001;
12'b100111111001: finv1 = 23'b00111011011010001001110;
12'b100111111010: finv1 = 23'b00111011010111000111100;
12'b100111111011: finv1 = 23'b00111011010100000101010;
12'b100111111100: finv1 = 23'b00111011010001000011001;
12'b100111111101: finv1 = 23'b00111011001110000001000;
12'b100111111110: finv1 = 23'b00111011001010111111000;
12'b100111111111: finv1 = 23'b00111011000111111101000;
12'b101000000000: finv1 = 23'b00111011000100111011001;
12'b101000000001: finv1 = 23'b00111011000001111001010;
12'b101000000010: finv1 = 23'b00111010111110110111011;
12'b101000000011: finv1 = 23'b00111010111011110101101;
12'b101000000100: finv1 = 23'b00111010111000110100000;
12'b101000000101: finv1 = 23'b00111010110101110010011;
12'b101000000110: finv1 = 23'b00111010110010110000110;
12'b101000000111: finv1 = 23'b00111010101111101111010;
12'b101000001000: finv1 = 23'b00111010101100101101110;
12'b101000001001: finv1 = 23'b00111010101001101100011;
12'b101000001010: finv1 = 23'b00111010100110101011000;
12'b101000001011: finv1 = 23'b00111010100011101001110;
12'b101000001100: finv1 = 23'b00111010100000101000100;
12'b101000001101: finv1 = 23'b00111010011101100111011;
12'b101000001110: finv1 = 23'b00111010011010100110010;
12'b101000001111: finv1 = 23'b00111010010111100101010;
12'b101000010000: finv1 = 23'b00111010010100100100010;
12'b101000010001: finv1 = 23'b00111010010001100011010;
12'b101000010010: finv1 = 23'b00111010001110100010011;
12'b101000010011: finv1 = 23'b00111010001011100001101;
12'b101000010100: finv1 = 23'b00111010001000100000111;
12'b101000010101: finv1 = 23'b00111010000101100000001;
12'b101000010110: finv1 = 23'b00111010000010011111100;
12'b101000010111: finv1 = 23'b00111001111111011110111;
12'b101000011000: finv1 = 23'b00111001111100011110011;
12'b101000011001: finv1 = 23'b00111001111001011101111;
12'b101000011010: finv1 = 23'b00111001110110011101100;
12'b101000011011: finv1 = 23'b00111001110011011101001;
12'b101000011100: finv1 = 23'b00111001110000011100110;
12'b101000011101: finv1 = 23'b00111001101101011100100;
12'b101000011110: finv1 = 23'b00111001101010011100011;
12'b101000011111: finv1 = 23'b00111001100111011100010;
12'b101000100000: finv1 = 23'b00111001100100011100001;
12'b101000100001: finv1 = 23'b00111001100001011100001;
12'b101000100010: finv1 = 23'b00111001011110011100010;
12'b101000100011: finv1 = 23'b00111001011011011100010;
12'b101000100100: finv1 = 23'b00111001011000011100100;
12'b101000100101: finv1 = 23'b00111001010101011100101;
12'b101000100110: finv1 = 23'b00111001010010011101000;
12'b101000100111: finv1 = 23'b00111001001111011101010;
12'b101000101000: finv1 = 23'b00111001001100011101101;
12'b101000101001: finv1 = 23'b00111001001001011110001;
12'b101000101010: finv1 = 23'b00111001000110011110101;
12'b101000101011: finv1 = 23'b00111001000011011111001;
12'b101000101100: finv1 = 23'b00111001000000011111110;
12'b101000101101: finv1 = 23'b00111000111101100000100;
12'b101000101110: finv1 = 23'b00111000111010100001010;
12'b101000101111: finv1 = 23'b00111000110111100010000;
12'b101000110000: finv1 = 23'b00111000110100100010111;
12'b101000110001: finv1 = 23'b00111000110001100011110;
12'b101000110010: finv1 = 23'b00111000101110100100101;
12'b101000110011: finv1 = 23'b00111000101011100101110;
12'b101000110100: finv1 = 23'b00111000101000100110110;
12'b101000110101: finv1 = 23'b00111000100101100111111;
12'b101000110110: finv1 = 23'b00111000100010101001001;
12'b101000110111: finv1 = 23'b00111000011111101010011;
12'b101000111000: finv1 = 23'b00111000011100101011101;
12'b101000111001: finv1 = 23'b00111000011001101101000;
12'b101000111010: finv1 = 23'b00111000010110101110011;
12'b101000111011: finv1 = 23'b00111000010011101111111;
12'b101000111100: finv1 = 23'b00111000010000110001011;
12'b101000111101: finv1 = 23'b00111000001101110011000;
12'b101000111110: finv1 = 23'b00111000001010110100101;
12'b101000111111: finv1 = 23'b00111000000111110110011;
12'b101001000000: finv1 = 23'b00111000000100111000001;
12'b101001000001: finv1 = 23'b00111000000001111001111;
12'b101001000010: finv1 = 23'b00110111111110111011110;
12'b101001000011: finv1 = 23'b00110111111011111101101;
12'b101001000100: finv1 = 23'b00110111111000111111101;
12'b101001000101: finv1 = 23'b00110111110110000001110;
12'b101001000110: finv1 = 23'b00110111110011000011110;
12'b101001000111: finv1 = 23'b00110111110000000101111;
12'b101001001000: finv1 = 23'b00110111101101001000001;
12'b101001001001: finv1 = 23'b00110111101010001010011;
12'b101001001010: finv1 = 23'b00110111100111001100110;
12'b101001001011: finv1 = 23'b00110111100100001111001;
12'b101001001100: finv1 = 23'b00110111100001010001100;
12'b101001001101: finv1 = 23'b00110111011110010100000;
12'b101001001110: finv1 = 23'b00110111011011010110101;
12'b101001001111: finv1 = 23'b00110111011000011001001;
12'b101001010000: finv1 = 23'b00110111010101011011111;
12'b101001010001: finv1 = 23'b00110111010010011110100;
12'b101001010010: finv1 = 23'b00110111001111100001010;
12'b101001010011: finv1 = 23'b00110111001100100100001;
12'b101001010100: finv1 = 23'b00110111001001100111000;
12'b101001010101: finv1 = 23'b00110111000110101010000;
12'b101001010110: finv1 = 23'b00110111000011101101000;
12'b101001010111: finv1 = 23'b00110111000000110000000;
12'b101001011000: finv1 = 23'b00110110111101110011001;
12'b101001011001: finv1 = 23'b00110110111010110110010;
12'b101001011010: finv1 = 23'b00110110110111111001100;
12'b101001011011: finv1 = 23'b00110110110100111100110;
12'b101001011100: finv1 = 23'b00110110110010000000001;
12'b101001011101: finv1 = 23'b00110110101111000011100;
12'b101001011110: finv1 = 23'b00110110101100000110111;
12'b101001011111: finv1 = 23'b00110110101001001010011;
12'b101001100000: finv1 = 23'b00110110100110001110000;
12'b101001100001: finv1 = 23'b00110110100011010001100;
12'b101001100010: finv1 = 23'b00110110100000010101010;
12'b101001100011: finv1 = 23'b00110110011101011001000;
12'b101001100100: finv1 = 23'b00110110011010011100110;
12'b101001100101: finv1 = 23'b00110110010111100000100;
12'b101001100110: finv1 = 23'b00110110010100100100100;
12'b101001100111: finv1 = 23'b00110110010001101000011;
12'b101001101000: finv1 = 23'b00110110001110101100011;
12'b101001101001: finv1 = 23'b00110110001011110000100;
12'b101001101010: finv1 = 23'b00110110001000110100100;
12'b101001101011: finv1 = 23'b00110110000101111000110;
12'b101001101100: finv1 = 23'b00110110000010111100111;
12'b101001101101: finv1 = 23'b00110110000000000001010;
12'b101001101110: finv1 = 23'b00110101111101000101100;
12'b101001101111: finv1 = 23'b00110101111010001001111;
12'b101001110000: finv1 = 23'b00110101110111001110011;
12'b101001110001: finv1 = 23'b00110101110100010010111;
12'b101001110010: finv1 = 23'b00110101110001010111011;
12'b101001110011: finv1 = 23'b00110101101110011100000;
12'b101001110100: finv1 = 23'b00110101101011100000110;
12'b101001110101: finv1 = 23'b00110101101000100101011;
12'b101001110110: finv1 = 23'b00110101100101101010010;
12'b101001110111: finv1 = 23'b00110101100010101111000;
12'b101001111000: finv1 = 23'b00110101011111110011111;
12'b101001111001: finv1 = 23'b00110101011100111000111;
12'b101001111010: finv1 = 23'b00110101011001111101111;
12'b101001111011: finv1 = 23'b00110101010111000010111;
12'b101001111100: finv1 = 23'b00110101010100001000000;
12'b101001111101: finv1 = 23'b00110101010001001101001;
12'b101001111110: finv1 = 23'b00110101001110010010011;
12'b101001111111: finv1 = 23'b00110101001011010111101;
12'b101010000000: finv1 = 23'b00110101001000011101000;
12'b101010000001: finv1 = 23'b00110101000101100010011;
12'b101010000010: finv1 = 23'b00110101000010100111110;
12'b101010000011: finv1 = 23'b00110100111111101101010;
12'b101010000100: finv1 = 23'b00110100111100110010111;
12'b101010000101: finv1 = 23'b00110100111001111000100;
12'b101010000110: finv1 = 23'b00110100110110111110001;
12'b101010000111: finv1 = 23'b00110100110100000011110;
12'b101010001000: finv1 = 23'b00110100110001001001101;
12'b101010001001: finv1 = 23'b00110100101110001111011;
12'b101010001010: finv1 = 23'b00110100101011010101010;
12'b101010001011: finv1 = 23'b00110100101000011011010;
12'b101010001100: finv1 = 23'b00110100100101100001001;
12'b101010001101: finv1 = 23'b00110100100010100111010;
12'b101010001110: finv1 = 23'b00110100011111101101011;
12'b101010001111: finv1 = 23'b00110100011100110011100;
12'b101010010000: finv1 = 23'b00110100011001111001101;
12'b101010010001: finv1 = 23'b00110100010110111111111;
12'b101010010010: finv1 = 23'b00110100010100000110010;
12'b101010010011: finv1 = 23'b00110100010001001100101;
12'b101010010100: finv1 = 23'b00110100001110010011000;
12'b101010010101: finv1 = 23'b00110100001011011001100;
12'b101010010110: finv1 = 23'b00110100001000100000000;
12'b101010010111: finv1 = 23'b00110100000101100110101;
12'b101010011000: finv1 = 23'b00110100000010101101010;
12'b101010011001: finv1 = 23'b00110011111111110100000;
12'b101010011010: finv1 = 23'b00110011111100111010110;
12'b101010011011: finv1 = 23'b00110011111010000001100;
12'b101010011100: finv1 = 23'b00110011110111001000011;
12'b101010011101: finv1 = 23'b00110011110100001111010;
12'b101010011110: finv1 = 23'b00110011110001010110010;
12'b101010011111: finv1 = 23'b00110011101110011101010;
12'b101010100000: finv1 = 23'b00110011101011100100011;
12'b101010100001: finv1 = 23'b00110011101000101011100;
12'b101010100010: finv1 = 23'b00110011100101110010101;
12'b101010100011: finv1 = 23'b00110011100010111001111;
12'b101010100100: finv1 = 23'b00110011100000000001010;
12'b101010100101: finv1 = 23'b00110011011101001000100;
12'b101010100110: finv1 = 23'b00110011011010010000000;
12'b101010100111: finv1 = 23'b00110011010111010111011;
12'b101010101000: finv1 = 23'b00110011010100011110111;
12'b101010101001: finv1 = 23'b00110011010001100110100;
12'b101010101010: finv1 = 23'b00110011001110101110001;
12'b101010101011: finv1 = 23'b00110011001011110101110;
12'b101010101100: finv1 = 23'b00110011001000111101100;
12'b101010101101: finv1 = 23'b00110011000110000101010;
12'b101010101110: finv1 = 23'b00110011000011001101001;
12'b101010101111: finv1 = 23'b00110011000000010101000;
12'b101010110000: finv1 = 23'b00110010111101011100111;
12'b101010110001: finv1 = 23'b00110010111010100100111;
12'b101010110010: finv1 = 23'b00110010110111101101000;
12'b101010110011: finv1 = 23'b00110010110100110101001;
12'b101010110100: finv1 = 23'b00110010110001111101010;
12'b101010110101: finv1 = 23'b00110010101111000101100;
12'b101010110110: finv1 = 23'b00110010101100001101110;
12'b101010110111: finv1 = 23'b00110010101001010110000;
12'b101010111000: finv1 = 23'b00110010100110011110011;
12'b101010111001: finv1 = 23'b00110010100011100110111;
12'b101010111010: finv1 = 23'b00110010100000101111010;
12'b101010111011: finv1 = 23'b00110010011101110111111;
12'b101010111100: finv1 = 23'b00110010011011000000011;
12'b101010111101: finv1 = 23'b00110010011000001001000;
12'b101010111110: finv1 = 23'b00110010010101010001110;
12'b101010111111: finv1 = 23'b00110010010010011010100;
12'b101011000000: finv1 = 23'b00110010001111100011010;
12'b101011000001: finv1 = 23'b00110010001100101100001;
12'b101011000010: finv1 = 23'b00110010001001110101000;
12'b101011000011: finv1 = 23'b00110010000110111110000;
12'b101011000100: finv1 = 23'b00110010000100000111000;
12'b101011000101: finv1 = 23'b00110010000001010000001;
12'b101011000110: finv1 = 23'b00110001111110011001010;
12'b101011000111: finv1 = 23'b00110001111011100010011;
12'b101011001000: finv1 = 23'b00110001111000101011101;
12'b101011001001: finv1 = 23'b00110001110101110100111;
12'b101011001010: finv1 = 23'b00110001110010111110010;
12'b101011001011: finv1 = 23'b00110001110000000111101;
12'b101011001100: finv1 = 23'b00110001101101010001000;
12'b101011001101: finv1 = 23'b00110001101010011010100;
12'b101011001110: finv1 = 23'b00110001100111100100001;
12'b101011001111: finv1 = 23'b00110001100100101101110;
12'b101011010000: finv1 = 23'b00110001100001110111011;
12'b101011010001: finv1 = 23'b00110001011111000001000;
12'b101011010010: finv1 = 23'b00110001011100001010111;
12'b101011010011: finv1 = 23'b00110001011001010100101;
12'b101011010100: finv1 = 23'b00110001010110011110100;
12'b101011010101: finv1 = 23'b00110001010011101000011;
12'b101011010110: finv1 = 23'b00110001010000110010011;
12'b101011010111: finv1 = 23'b00110001001101111100011;
12'b101011011000: finv1 = 23'b00110001001011000110100;
12'b101011011001: finv1 = 23'b00110001001000010000101;
12'b101011011010: finv1 = 23'b00110001000101011010110;
12'b101011011011: finv1 = 23'b00110001000010100101000;
12'b101011011100: finv1 = 23'b00110000111111101111011;
12'b101011011101: finv1 = 23'b00110000111100111001101;
12'b101011011110: finv1 = 23'b00110000111010000100000;
12'b101011011111: finv1 = 23'b00110000110111001110100;
12'b101011100000: finv1 = 23'b00110000110100011001000;
12'b101011100001: finv1 = 23'b00110000110001100011100;
12'b101011100010: finv1 = 23'b00110000101110101110001;
12'b101011100011: finv1 = 23'b00110000101011111000111;
12'b101011100100: finv1 = 23'b00110000101001000011100;
12'b101011100101: finv1 = 23'b00110000100110001110010;
12'b101011100110: finv1 = 23'b00110000100011011001001;
12'b101011100111: finv1 = 23'b00110000100000100100000;
12'b101011101000: finv1 = 23'b00110000011101101110111;
12'b101011101001: finv1 = 23'b00110000011010111001111;
12'b101011101010: finv1 = 23'b00110000011000000100111;
12'b101011101011: finv1 = 23'b00110000010101010000000;
12'b101011101100: finv1 = 23'b00110000010010011011001;
12'b101011101101: finv1 = 23'b00110000001111100110010;
12'b101011101110: finv1 = 23'b00110000001100110001100;
12'b101011101111: finv1 = 23'b00110000001001111100111;
12'b101011110000: finv1 = 23'b00110000000111001000001;
12'b101011110001: finv1 = 23'b00110000000100010011100;
12'b101011110010: finv1 = 23'b00110000000001011111000;
12'b101011110011: finv1 = 23'b00101111111110101010100;
12'b101011110100: finv1 = 23'b00101111111011110110000;
12'b101011110101: finv1 = 23'b00101111111001000001101;
12'b101011110110: finv1 = 23'b00101111110110001101011;
12'b101011110111: finv1 = 23'b00101111110011011001000;
12'b101011111000: finv1 = 23'b00101111110000100100110;
12'b101011111001: finv1 = 23'b00101111101101110000101;
12'b101011111010: finv1 = 23'b00101111101010111100100;
12'b101011111011: finv1 = 23'b00101111101000001000011;
12'b101011111100: finv1 = 23'b00101111100101010100011;
12'b101011111101: finv1 = 23'b00101111100010100000011;
12'b101011111110: finv1 = 23'b00101111011111101100100;
12'b101011111111: finv1 = 23'b00101111011100111000101;
12'b101100000000: finv1 = 23'b00101111011010000100110;
12'b101100000001: finv1 = 23'b00101111010111010001000;
12'b101100000010: finv1 = 23'b00101111010100011101010;
12'b101100000011: finv1 = 23'b00101111010001101001101;
12'b101100000100: finv1 = 23'b00101111001110110110000;
12'b101100000101: finv1 = 23'b00101111001100000010011;
12'b101100000110: finv1 = 23'b00101111001001001110111;
12'b101100000111: finv1 = 23'b00101111000110011011011;
12'b101100001000: finv1 = 23'b00101111000011101000000;
12'b101100001001: finv1 = 23'b00101111000000110100101;
12'b101100001010: finv1 = 23'b00101110111110000001011;
12'b101100001011: finv1 = 23'b00101110111011001110001;
12'b101100001100: finv1 = 23'b00101110111000011010111;
12'b101100001101: finv1 = 23'b00101110110101100111110;
12'b101100001110: finv1 = 23'b00101110110010110100101;
12'b101100001111: finv1 = 23'b00101110110000000001101;
12'b101100010000: finv1 = 23'b00101110101101001110101;
12'b101100010001: finv1 = 23'b00101110101010011011110;
12'b101100010010: finv1 = 23'b00101110100111101000110;
12'b101100010011: finv1 = 23'b00101110100100110110000;
12'b101100010100: finv1 = 23'b00101110100010000011001;
12'b101100010101: finv1 = 23'b00101110011111010000100;
12'b101100010110: finv1 = 23'b00101110011100011101110;
12'b101100010111: finv1 = 23'b00101110011001101011001;
12'b101100011000: finv1 = 23'b00101110010110111000100;
12'b101100011001: finv1 = 23'b00101110010100000110000;
12'b101100011010: finv1 = 23'b00101110010001010011100;
12'b101100011011: finv1 = 23'b00101110001110100001001;
12'b101100011100: finv1 = 23'b00101110001011101110110;
12'b101100011101: finv1 = 23'b00101110001000111100011;
12'b101100011110: finv1 = 23'b00101110000110001010001;
12'b101100011111: finv1 = 23'b00101110000011010111111;
12'b101100100000: finv1 = 23'b00101110000000100101110;
12'b101100100001: finv1 = 23'b00101101111101110011101;
12'b101100100010: finv1 = 23'b00101101111011000001101;
12'b101100100011: finv1 = 23'b00101101111000001111100;
12'b101100100100: finv1 = 23'b00101101110101011101101;
12'b101100100101: finv1 = 23'b00101101110010101011101;
12'b101100100110: finv1 = 23'b00101101101111111001110;
12'b101100100111: finv1 = 23'b00101101101101001000000;
12'b101100101000: finv1 = 23'b00101101101010010110010;
12'b101100101001: finv1 = 23'b00101101100111100100100;
12'b101100101010: finv1 = 23'b00101101100100110010111;
12'b101100101011: finv1 = 23'b00101101100010000001010;
12'b101100101100: finv1 = 23'b00101101011111001111110;
12'b101100101101: finv1 = 23'b00101101011100011110010;
12'b101100101110: finv1 = 23'b00101101011001101100110;
12'b101100101111: finv1 = 23'b00101101010110111011011;
12'b101100110000: finv1 = 23'b00101101010100001010000;
12'b101100110001: finv1 = 23'b00101101010001011000110;
12'b101100110010: finv1 = 23'b00101101001110100111100;
12'b101100110011: finv1 = 23'b00101101001011110110010;
12'b101100110100: finv1 = 23'b00101101001001000101001;
12'b101100110101: finv1 = 23'b00101101000110010100000;
12'b101100110110: finv1 = 23'b00101101000011100011000;
12'b101100110111: finv1 = 23'b00101101000000110010000;
12'b101100111000: finv1 = 23'b00101100111110000001000;
12'b101100111001: finv1 = 23'b00101100111011010000001;
12'b101100111010: finv1 = 23'b00101100111000011111010;
12'b101100111011: finv1 = 23'b00101100110101101110100;
12'b101100111100: finv1 = 23'b00101100110010111101110;
12'b101100111101: finv1 = 23'b00101100110000001101001;
12'b101100111110: finv1 = 23'b00101100101101011100011;
12'b101100111111: finv1 = 23'b00101100101010101011111;
12'b101101000000: finv1 = 23'b00101100100111111011010;
12'b101101000001: finv1 = 23'b00101100100101001010111;
12'b101101000010: finv1 = 23'b00101100100010011010011;
12'b101101000011: finv1 = 23'b00101100011111101010000;
12'b101101000100: finv1 = 23'b00101100011100111001101;
12'b101101000101: finv1 = 23'b00101100011010001001011;
12'b101101000110: finv1 = 23'b00101100010111011001001;
12'b101101000111: finv1 = 23'b00101100010100101001000;
12'b101101001000: finv1 = 23'b00101100010001111000111;
12'b101101001001: finv1 = 23'b00101100001111001000110;
12'b101101001010: finv1 = 23'b00101100001100011000110;
12'b101101001011: finv1 = 23'b00101100001001101000110;
12'b101101001100: finv1 = 23'b00101100000110111000110;
12'b101101001101: finv1 = 23'b00101100000100001000111;
12'b101101001110: finv1 = 23'b00101100000001011001001;
12'b101101001111: finv1 = 23'b00101011111110101001010;
12'b101101010000: finv1 = 23'b00101011111011111001100;
12'b101101010001: finv1 = 23'b00101011111001001001111;
12'b101101010010: finv1 = 23'b00101011110110011010010;
12'b101101010011: finv1 = 23'b00101011110011101010101;
12'b101101010100: finv1 = 23'b00101011110000111011001;
12'b101101010101: finv1 = 23'b00101011101110001011101;
12'b101101010110: finv1 = 23'b00101011101011011100010;
12'b101101010111: finv1 = 23'b00101011101000101100111;
12'b101101011000: finv1 = 23'b00101011100101111101100;
12'b101101011001: finv1 = 23'b00101011100011001110010;
12'b101101011010: finv1 = 23'b00101011100000011111000;
12'b101101011011: finv1 = 23'b00101011011101101111111;
12'b101101011100: finv1 = 23'b00101011011011000000110;
12'b101101011101: finv1 = 23'b00101011011000010001101;
12'b101101011110: finv1 = 23'b00101011010101100010101;
12'b101101011111: finv1 = 23'b00101011010010110011101;
12'b101101100000: finv1 = 23'b00101011010000000100101;
12'b101101100001: finv1 = 23'b00101011001101010101110;
12'b101101100010: finv1 = 23'b00101011001010100111000;
12'b101101100011: finv1 = 23'b00101011000111111000001;
12'b101101100100: finv1 = 23'b00101011000101001001100;
12'b101101100101: finv1 = 23'b00101011000010011010110;
12'b101101100110: finv1 = 23'b00101010111111101100001;
12'b101101100111: finv1 = 23'b00101010111100111101101;
12'b101101101000: finv1 = 23'b00101010111010001111000;
12'b101101101001: finv1 = 23'b00101010110111100000100;
12'b101101101010: finv1 = 23'b00101010110100110010001;
12'b101101101011: finv1 = 23'b00101010110010000011110;
12'b101101101100: finv1 = 23'b00101010101111010101011;
12'b101101101101: finv1 = 23'b00101010101100100111001;
12'b101101101110: finv1 = 23'b00101010101001111000111;
12'b101101101111: finv1 = 23'b00101010100111001010110;
12'b101101110000: finv1 = 23'b00101010100100011100101;
12'b101101110001: finv1 = 23'b00101010100001101110100;
12'b101101110010: finv1 = 23'b00101010011111000000100;
12'b101101110011: finv1 = 23'b00101010011100010010100;
12'b101101110100: finv1 = 23'b00101010011001100100100;
12'b101101110101: finv1 = 23'b00101010010110110110101;
12'b101101110110: finv1 = 23'b00101010010100001000111;
12'b101101110111: finv1 = 23'b00101010010001011011000;
12'b101101111000: finv1 = 23'b00101010001110101101010;
12'b101101111001: finv1 = 23'b00101010001011111111101;
12'b101101111010: finv1 = 23'b00101010001001010010000;
12'b101101111011: finv1 = 23'b00101010000110100100011;
12'b101101111100: finv1 = 23'b00101010000011110110111;
12'b101101111101: finv1 = 23'b00101010000001001001011;
12'b101101111110: finv1 = 23'b00101001111110011011111;
12'b101101111111: finv1 = 23'b00101001111011101110100;
12'b101110000000: finv1 = 23'b00101001111001000001001;
12'b101110000001: finv1 = 23'b00101001110110010011111;
12'b101110000010: finv1 = 23'b00101001110011100110101;
12'b101110000011: finv1 = 23'b00101001110000111001011;
12'b101110000100: finv1 = 23'b00101001101110001100010;
12'b101110000101: finv1 = 23'b00101001101011011111001;
12'b101110000110: finv1 = 23'b00101001101000110010001;
12'b101110000111: finv1 = 23'b00101001100110000101001;
12'b101110001000: finv1 = 23'b00101001100011011000010;
12'b101110001001: finv1 = 23'b00101001100000101011010;
12'b101110001010: finv1 = 23'b00101001011101111110100;
12'b101110001011: finv1 = 23'b00101001011011010001101;
12'b101110001100: finv1 = 23'b00101001011000100100111;
12'b101110001101: finv1 = 23'b00101001010101111000001;
12'b101110001110: finv1 = 23'b00101001010011001011100;
12'b101110001111: finv1 = 23'b00101001010000011110111;
12'b101110010000: finv1 = 23'b00101001001101110010011;
12'b101110010001: finv1 = 23'b00101001001011000101111;
12'b101110010010: finv1 = 23'b00101001001000011001011;
12'b101110010011: finv1 = 23'b00101001000101101101000;
12'b101110010100: finv1 = 23'b00101001000011000000101;
12'b101110010101: finv1 = 23'b00101001000000010100010;
12'b101110010110: finv1 = 23'b00101000111101101000000;
12'b101110010111: finv1 = 23'b00101000111010111011111;
12'b101110011000: finv1 = 23'b00101000111000001111101;
12'b101110011001: finv1 = 23'b00101000110101100011100;
12'b101110011010: finv1 = 23'b00101000110010110111100;
12'b101110011011: finv1 = 23'b00101000110000001011100;
12'b101110011100: finv1 = 23'b00101000101101011111100;
12'b101110011101: finv1 = 23'b00101000101010110011100;
12'b101110011110: finv1 = 23'b00101000101000000111101;
12'b101110011111: finv1 = 23'b00101000100101011011111;
12'b101110100000: finv1 = 23'b00101000100010110000001;
12'b101110100001: finv1 = 23'b00101000100000000100011;
12'b101110100010: finv1 = 23'b00101000011101011000101;
12'b101110100011: finv1 = 23'b00101000011010101101000;
12'b101110100100: finv1 = 23'b00101000011000000001100;
12'b101110100101: finv1 = 23'b00101000010101010101111;
12'b101110100110: finv1 = 23'b00101000010010101010011;
12'b101110100111: finv1 = 23'b00101000001111111111000;
12'b101110101000: finv1 = 23'b00101000001101010011101;
12'b101110101001: finv1 = 23'b00101000001010101000010;
12'b101110101010: finv1 = 23'b00101000000111111101000;
12'b101110101011: finv1 = 23'b00101000000101010001110;
12'b101110101100: finv1 = 23'b00101000000010100110100;
12'b101110101101: finv1 = 23'b00100111111111111011011;
12'b101110101110: finv1 = 23'b00100111111101010000010;
12'b101110101111: finv1 = 23'b00100111111010100101010;
12'b101110110000: finv1 = 23'b00100111110111111010010;
12'b101110110001: finv1 = 23'b00100111110101001111010;
12'b101110110010: finv1 = 23'b00100111110010100100011;
12'b101110110011: finv1 = 23'b00100111101111111001100;
12'b101110110100: finv1 = 23'b00100111101101001110110;
12'b101110110101: finv1 = 23'b00100111101010100011111;
12'b101110110110: finv1 = 23'b00100111100111111001010;
12'b101110110111: finv1 = 23'b00100111100101001110100;
12'b101110111000: finv1 = 23'b00100111100010100011111;
12'b101110111001: finv1 = 23'b00100111011111111001011;
12'b101110111010: finv1 = 23'b00100111011101001110111;
12'b101110111011: finv1 = 23'b00100111011010100100011;
12'b101110111100: finv1 = 23'b00100111010111111010000;
12'b101110111101: finv1 = 23'b00100111010101001111101;
12'b101110111110: finv1 = 23'b00100111010010100101010;
12'b101110111111: finv1 = 23'b00100111001111111011000;
12'b101111000000: finv1 = 23'b00100111001101010000110;
12'b101111000001: finv1 = 23'b00100111001010100110100;
12'b101111000010: finv1 = 23'b00100111000111111100011;
12'b101111000011: finv1 = 23'b00100111000101010010010;
12'b101111000100: finv1 = 23'b00100111000010101000010;
12'b101111000101: finv1 = 23'b00100110111111111110010;
12'b101111000110: finv1 = 23'b00100110111101010100011;
12'b101111000111: finv1 = 23'b00100110111010101010011;
12'b101111001000: finv1 = 23'b00100110111000000000101;
12'b101111001001: finv1 = 23'b00100110110101010110110;
12'b101111001010: finv1 = 23'b00100110110010101101000;
12'b101111001011: finv1 = 23'b00100110110000000011010;
12'b101111001100: finv1 = 23'b00100110101101011001101;
12'b101111001101: finv1 = 23'b00100110101010110000000;
12'b101111001110: finv1 = 23'b00100110101000000110100;
12'b101111001111: finv1 = 23'b00100110100101011101000;
12'b101111010000: finv1 = 23'b00100110100010110011100;
12'b101111010001: finv1 = 23'b00100110100000001010001;
12'b101111010010: finv1 = 23'b00100110011101100000110;
12'b101111010011: finv1 = 23'b00100110011010110111011;
12'b101111010100: finv1 = 23'b00100110011000001110001;
12'b101111010101: finv1 = 23'b00100110010101100100111;
12'b101111010110: finv1 = 23'b00100110010010111011101;
12'b101111010111: finv1 = 23'b00100110010000010010100;
12'b101111011000: finv1 = 23'b00100110001101101001100;
12'b101111011001: finv1 = 23'b00100110001011000000011;
12'b101111011010: finv1 = 23'b00100110001000010111011;
12'b101111011011: finv1 = 23'b00100110000101101110100;
12'b101111011100: finv1 = 23'b00100110000011000101101;
12'b101111011101: finv1 = 23'b00100110000000011100110;
12'b101111011110: finv1 = 23'b00100101111101110011111;
12'b101111011111: finv1 = 23'b00100101111011001011001;
12'b101111100000: finv1 = 23'b00100101111000100010100;
12'b101111100001: finv1 = 23'b00100101110101111001110;
12'b101111100010: finv1 = 23'b00100101110011010001001;
12'b101111100011: finv1 = 23'b00100101110000101000101;
12'b101111100100: finv1 = 23'b00100101101110000000001;
12'b101111100101: finv1 = 23'b00100101101011010111101;
12'b101111100110: finv1 = 23'b00100101101000101111001;
12'b101111100111: finv1 = 23'b00100101100110000110110;
12'b101111101000: finv1 = 23'b00100101100011011110100;
12'b101111101001: finv1 = 23'b00100101100000110110001;
12'b101111101010: finv1 = 23'b00100101011110001101111;
12'b101111101011: finv1 = 23'b00100101011011100101110;
12'b101111101100: finv1 = 23'b00100101011000111101101;
12'b101111101101: finv1 = 23'b00100101010110010101100;
12'b101111101110: finv1 = 23'b00100101010011101101100;
12'b101111101111: finv1 = 23'b00100101010001000101100;
12'b101111110000: finv1 = 23'b00100101001110011101100;
12'b101111110001: finv1 = 23'b00100101001011110101101;
12'b101111110010: finv1 = 23'b00100101001001001101110;
12'b101111110011: finv1 = 23'b00100101000110100101111;
12'b101111110100: finv1 = 23'b00100101000011111110001;
12'b101111110101: finv1 = 23'b00100101000001010110011;
12'b101111110110: finv1 = 23'b00100100111110101110110;
12'b101111110111: finv1 = 23'b00100100111100000111001;
12'b101111111000: finv1 = 23'b00100100111001011111100;
12'b101111111001: finv1 = 23'b00100100110110111000000;
12'b101111111010: finv1 = 23'b00100100110100010000100;
12'b101111111011: finv1 = 23'b00100100110001101001001;
12'b101111111100: finv1 = 23'b00100100101111000001101;
12'b101111111101: finv1 = 23'b00100100101100011010011;
12'b101111111110: finv1 = 23'b00100100101001110011000;
12'b101111111111: finv1 = 23'b00100100100111001011110;
12'b110000000000: finv1 = 23'b00100100100100100100101;
12'b110000000001: finv1 = 23'b00100100100001111101011;
12'b110000000010: finv1 = 23'b00100100011111010110010;
12'b110000000011: finv1 = 23'b00100100011100101111010;
12'b110000000100: finv1 = 23'b00100100011010001000010;
12'b110000000101: finv1 = 23'b00100100010111100001010;
12'b110000000110: finv1 = 23'b00100100010100111010010;
12'b110000000111: finv1 = 23'b00100100010010010011011;
12'b110000001000: finv1 = 23'b00100100001111101100101;
12'b110000001001: finv1 = 23'b00100100001101000101110;
12'b110000001010: finv1 = 23'b00100100001010011111001;
12'b110000001011: finv1 = 23'b00100100000111111000011;
12'b110000001100: finv1 = 23'b00100100000101010001110;
12'b110000001101: finv1 = 23'b00100100000010101011001;
12'b110000001110: finv1 = 23'b00100100000000000100101;
12'b110000001111: finv1 = 23'b00100011111101011110000;
12'b110000010000: finv1 = 23'b00100011111010110111101;
12'b110000010001: finv1 = 23'b00100011111000010001001;
12'b110000010010: finv1 = 23'b00100011110101101010110;
12'b110000010011: finv1 = 23'b00100011110011000100100;
12'b110000010100: finv1 = 23'b00100011110000011110010;
12'b110000010101: finv1 = 23'b00100011101101111000000;
12'b110000010110: finv1 = 23'b00100011101011010001110;
12'b110000010111: finv1 = 23'b00100011101000101011101;
12'b110000011000: finv1 = 23'b00100011100110000101100;
12'b110000011001: finv1 = 23'b00100011100011011111100;
12'b110000011010: finv1 = 23'b00100011100000111001100;
12'b110000011011: finv1 = 23'b00100011011110010011100;
12'b110000011100: finv1 = 23'b00100011011011101101101;
12'b110000011101: finv1 = 23'b00100011011001000111110;
12'b110000011110: finv1 = 23'b00100011010110100010000;
12'b110000011111: finv1 = 23'b00100011010011111100010;
12'b110000100000: finv1 = 23'b00100011010001010110100;
12'b110000100001: finv1 = 23'b00100011001110110000110;
12'b110000100010: finv1 = 23'b00100011001100001011001;
12'b110000100011: finv1 = 23'b00100011001001100101101;
12'b110000100100: finv1 = 23'b00100011000111000000000;
12'b110000100101: finv1 = 23'b00100011000100011010100;
12'b110000100110: finv1 = 23'b00100011000001110101001;
12'b110000100111: finv1 = 23'b00100010111111001111110;
12'b110000101000: finv1 = 23'b00100010111100101010011;
12'b110000101001: finv1 = 23'b00100010111010000101000;
12'b110000101010: finv1 = 23'b00100010110111011111110;
12'b110000101011: finv1 = 23'b00100010110100111010100;
12'b110000101100: finv1 = 23'b00100010110010010101011;
12'b110000101101: finv1 = 23'b00100010101111110000010;
12'b110000101110: finv1 = 23'b00100010101101001011001;
12'b110000101111: finv1 = 23'b00100010101010100110001;
12'b110000110000: finv1 = 23'b00100010101000000001001;
12'b110000110001: finv1 = 23'b00100010100101011100010;
12'b110000110010: finv1 = 23'b00100010100010110111010;
12'b110000110011: finv1 = 23'b00100010100000010010100;
12'b110000110100: finv1 = 23'b00100010011101101101101;
12'b110000110101: finv1 = 23'b00100010011011001000111;
12'b110000110110: finv1 = 23'b00100010011000100100001;
12'b110000110111: finv1 = 23'b00100010010101111111100;
12'b110000111000: finv1 = 23'b00100010010011011010111;
12'b110000111001: finv1 = 23'b00100010010000110110010;
12'b110000111010: finv1 = 23'b00100010001110010001110;
12'b110000111011: finv1 = 23'b00100010001011101101010;
12'b110000111100: finv1 = 23'b00100010001001001000111;
12'b110000111101: finv1 = 23'b00100010000110100100011;
12'b110000111110: finv1 = 23'b00100010000100000000001;
12'b110000111111: finv1 = 23'b00100010000001011011110;
12'b110001000000: finv1 = 23'b00100001111110110111100;
12'b110001000001: finv1 = 23'b00100001111100010011010;
12'b110001000010: finv1 = 23'b00100001111001101111001;
12'b110001000011: finv1 = 23'b00100001110111001011000;
12'b110001000100: finv1 = 23'b00100001110100100110111;
12'b110001000101: finv1 = 23'b00100001110010000010111;
12'b110001000110: finv1 = 23'b00100001101111011110111;
12'b110001000111: finv1 = 23'b00100001101100111011000;
12'b110001001000: finv1 = 23'b00100001101010010111000;
12'b110001001001: finv1 = 23'b00100001100111110011010;
12'b110001001010: finv1 = 23'b00100001100101001111011;
12'b110001001011: finv1 = 23'b00100001100010101011101;
12'b110001001100: finv1 = 23'b00100001100000000111111;
12'b110001001101: finv1 = 23'b00100001011101100100010;
12'b110001001110: finv1 = 23'b00100001011011000000101;
12'b110001001111: finv1 = 23'b00100001011000011101000;
12'b110001010000: finv1 = 23'b00100001010101111001100;
12'b110001010001: finv1 = 23'b00100001010011010110000;
12'b110001010010: finv1 = 23'b00100001010000110010101;
12'b110001010011: finv1 = 23'b00100001001110001111001;
12'b110001010100: finv1 = 23'b00100001001011101011110;
12'b110001010101: finv1 = 23'b00100001001001001000100;
12'b110001010110: finv1 = 23'b00100001000110100101010;
12'b110001010111: finv1 = 23'b00100001000100000010000;
12'b110001011000: finv1 = 23'b00100001000001011110111;
12'b110001011001: finv1 = 23'b00100000111110111011110;
12'b110001011010: finv1 = 23'b00100000111100011000101;
12'b110001011011: finv1 = 23'b00100000111001110101101;
12'b110001011100: finv1 = 23'b00100000110111010010101;
12'b110001011101: finv1 = 23'b00100000110100101111101;
12'b110001011110: finv1 = 23'b00100000110010001100110;
12'b110001011111: finv1 = 23'b00100000101111101001111;
12'b110001100000: finv1 = 23'b00100000101101000111000;
12'b110001100001: finv1 = 23'b00100000101010100100010;
12'b110001100010: finv1 = 23'b00100000101000000001100;
12'b110001100011: finv1 = 23'b00100000100101011110111;
12'b110001100100: finv1 = 23'b00100000100010111100010;
12'b110001100101: finv1 = 23'b00100000100000011001101;
12'b110001100110: finv1 = 23'b00100000011101110111001;
12'b110001100111: finv1 = 23'b00100000011011010100101;
12'b110001101000: finv1 = 23'b00100000011000110010001;
12'b110001101001: finv1 = 23'b00100000010110001111110;
12'b110001101010: finv1 = 23'b00100000010011101101011;
12'b110001101011: finv1 = 23'b00100000010001001011000;
12'b110001101100: finv1 = 23'b00100000001110101000110;
12'b110001101101: finv1 = 23'b00100000001100000110100;
12'b110001101110: finv1 = 23'b00100000001001100100011;
12'b110001101111: finv1 = 23'b00100000000111000010001;
12'b110001110000: finv1 = 23'b00100000000100100000001;
12'b110001110001: finv1 = 23'b00100000000001111110000;
12'b110001110010: finv1 = 23'b00011111111111011100000;
12'b110001110011: finv1 = 23'b00011111111100111010000;
12'b110001110100: finv1 = 23'b00011111111010011000001;
12'b110001110101: finv1 = 23'b00011111110111110110010;
12'b110001110110: finv1 = 23'b00011111110101010100011;
12'b110001110111: finv1 = 23'b00011111110010110010101;
12'b110001111000: finv1 = 23'b00011111110000010000111;
12'b110001111001: finv1 = 23'b00011111101101101111001;
12'b110001111010: finv1 = 23'b00011111101011001101100;
12'b110001111011: finv1 = 23'b00011111101000101011111;
12'b110001111100: finv1 = 23'b00011111100110001010011;
12'b110001111101: finv1 = 23'b00011111100011101000110;
12'b110001111110: finv1 = 23'b00011111100001000111011;
12'b110001111111: finv1 = 23'b00011111011110100101111;
12'b110010000000: finv1 = 23'b00011111011100000100100;
12'b110010000001: finv1 = 23'b00011111011001100011001;
12'b110010000010: finv1 = 23'b00011111010111000001111;
12'b110010000011: finv1 = 23'b00011111010100100000101;
12'b110010000100: finv1 = 23'b00011111010001111111011;
12'b110010000101: finv1 = 23'b00011111001111011110010;
12'b110010000110: finv1 = 23'b00011111001100111101001;
12'b110010000111: finv1 = 23'b00011111001010011100000;
12'b110010001000: finv1 = 23'b00011111000111111011000;
12'b110010001001: finv1 = 23'b00011111000101011010000;
12'b110010001010: finv1 = 23'b00011111000010111001000;
12'b110010001011: finv1 = 23'b00011111000000011000001;
12'b110010001100: finv1 = 23'b00011110111101110111010;
12'b110010001101: finv1 = 23'b00011110111011010110011;
12'b110010001110: finv1 = 23'b00011110111000110101101;
12'b110010001111: finv1 = 23'b00011110110110010100111;
12'b110010010000: finv1 = 23'b00011110110011110100010;
12'b110010010001: finv1 = 23'b00011110110001010011101;
12'b110010010010: finv1 = 23'b00011110101110110011000;
12'b110010010011: finv1 = 23'b00011110101100010010100;
12'b110010010100: finv1 = 23'b00011110101001110001111;
12'b110010010101: finv1 = 23'b00011110100111010001100;
12'b110010010110: finv1 = 23'b00011110100100110001000;
12'b110010010111: finv1 = 23'b00011110100010010000101;
12'b110010011000: finv1 = 23'b00011110011111110000011;
12'b110010011001: finv1 = 23'b00011110011101010000000;
12'b110010011010: finv1 = 23'b00011110011010101111110;
12'b110010011011: finv1 = 23'b00011110011000001111101;
12'b110010011100: finv1 = 23'b00011110010101101111011;
12'b110010011101: finv1 = 23'b00011110010011001111011;
12'b110010011110: finv1 = 23'b00011110010000101111010;
12'b110010011111: finv1 = 23'b00011110001110001111010;
12'b110010100000: finv1 = 23'b00011110001011101111010;
12'b110010100001: finv1 = 23'b00011110001001001111010;
12'b110010100010: finv1 = 23'b00011110000110101111011;
12'b110010100011: finv1 = 23'b00011110000100001111100;
12'b110010100100: finv1 = 23'b00011110000001101111110;
12'b110010100101: finv1 = 23'b00011101111111010000000;
12'b110010100110: finv1 = 23'b00011101111100110000010;
12'b110010100111: finv1 = 23'b00011101111010010000100;
12'b110010101000: finv1 = 23'b00011101110111110000111;
12'b110010101001: finv1 = 23'b00011101110101010001011;
12'b110010101010: finv1 = 23'b00011101110010110001110;
12'b110010101011: finv1 = 23'b00011101110000010010010;
12'b110010101100: finv1 = 23'b00011101101101110010111;
12'b110010101101: finv1 = 23'b00011101101011010011011;
12'b110010101110: finv1 = 23'b00011101101000110100000;
12'b110010101111: finv1 = 23'b00011101100110010100110;
12'b110010110000: finv1 = 23'b00011101100011110101011;
12'b110010110001: finv1 = 23'b00011101100001010110001;
12'b110010110010: finv1 = 23'b00011101011110110111000;
12'b110010110011: finv1 = 23'b00011101011100010111110;
12'b110010110100: finv1 = 23'b00011101011001111000101;
12'b110010110101: finv1 = 23'b00011101010111011001101;
12'b110010110110: finv1 = 23'b00011101010100111010101;
12'b110010110111: finv1 = 23'b00011101010010011011101;
12'b110010111000: finv1 = 23'b00011101001111111100101;
12'b110010111001: finv1 = 23'b00011101001101011101110;
12'b110010111010: finv1 = 23'b00011101001010111110111;
12'b110010111011: finv1 = 23'b00011101001000100000001;
12'b110010111100: finv1 = 23'b00011101000110000001011;
12'b110010111101: finv1 = 23'b00011101000011100010101;
12'b110010111110: finv1 = 23'b00011101000001000011111;
12'b110010111111: finv1 = 23'b00011100111110100101010;
12'b110011000000: finv1 = 23'b00011100111100000110101;
12'b110011000001: finv1 = 23'b00011100111001101000001;
12'b110011000010: finv1 = 23'b00011100110111001001101;
12'b110011000011: finv1 = 23'b00011100110100101011001;
12'b110011000100: finv1 = 23'b00011100110010001100110;
12'b110011000101: finv1 = 23'b00011100101111101110011;
12'b110011000110: finv1 = 23'b00011100101101010000000;
12'b110011000111: finv1 = 23'b00011100101010110001110;
12'b110011001000: finv1 = 23'b00011100101000010011100;
12'b110011001001: finv1 = 23'b00011100100101110101010;
12'b110011001010: finv1 = 23'b00011100100011010111001;
12'b110011001011: finv1 = 23'b00011100100000111001000;
12'b110011001100: finv1 = 23'b00011100011110011010111;
12'b110011001101: finv1 = 23'b00011100011011111100111;
12'b110011001110: finv1 = 23'b00011100011001011110111;
12'b110011001111: finv1 = 23'b00011100010111000000111;
12'b110011010000: finv1 = 23'b00011100010100100011000;
12'b110011010001: finv1 = 23'b00011100010010000101001;
12'b110011010010: finv1 = 23'b00011100001111100111010;
12'b110011010011: finv1 = 23'b00011100001101001001100;
12'b110011010100: finv1 = 23'b00011100001010101011110;
12'b110011010101: finv1 = 23'b00011100001000001110001;
12'b110011010110: finv1 = 23'b00011100000101110000011;
12'b110011010111: finv1 = 23'b00011100000011010010111;
12'b110011011000: finv1 = 23'b00011100000000110101010;
12'b110011011001: finv1 = 23'b00011011111110010111110;
12'b110011011010: finv1 = 23'b00011011111011111010010;
12'b110011011011: finv1 = 23'b00011011111001011100110;
12'b110011011100: finv1 = 23'b00011011110110111111011;
12'b110011011101: finv1 = 23'b00011011110100100010000;
12'b110011011110: finv1 = 23'b00011011110010000100110;
12'b110011011111: finv1 = 23'b00011011101111100111100;
12'b110011100000: finv1 = 23'b00011011101101001010010;
12'b110011100001: finv1 = 23'b00011011101010101101001;
12'b110011100010: finv1 = 23'b00011011101000001111111;
12'b110011100011: finv1 = 23'b00011011100101110010111;
12'b110011100100: finv1 = 23'b00011011100011010101110;
12'b110011100101: finv1 = 23'b00011011100000111000110;
12'b110011100110: finv1 = 23'b00011011011110011011110;
12'b110011100111: finv1 = 23'b00011011011011111110111;
12'b110011101000: finv1 = 23'b00011011011001100010000;
12'b110011101001: finv1 = 23'b00011011010111000101001;
12'b110011101010: finv1 = 23'b00011011010100101000011;
12'b110011101011: finv1 = 23'b00011011010010001011101;
12'b110011101100: finv1 = 23'b00011011001111101110111;
12'b110011101101: finv1 = 23'b00011011001101010010001;
12'b110011101110: finv1 = 23'b00011011001010110101100;
12'b110011101111: finv1 = 23'b00011011001000011001000;
12'b110011110000: finv1 = 23'b00011011000101111100011;
12'b110011110001: finv1 = 23'b00011011000011011111111;
12'b110011110010: finv1 = 23'b00011011000001000011100;
12'b110011110011: finv1 = 23'b00011010111110100111000;
12'b110011110100: finv1 = 23'b00011010111100001010101;
12'b110011110101: finv1 = 23'b00011010111001101110010;
12'b110011110110: finv1 = 23'b00011010110111010010000;
12'b110011110111: finv1 = 23'b00011010110100110101110;
12'b110011111000: finv1 = 23'b00011010110010011001100;
12'b110011111001: finv1 = 23'b00011010101111111101011;
12'b110011111010: finv1 = 23'b00011010101101100001010;
12'b110011111011: finv1 = 23'b00011010101011000101001;
12'b110011111100: finv1 = 23'b00011010101000101001001;
12'b110011111101: finv1 = 23'b00011010100110001101001;
12'b110011111110: finv1 = 23'b00011010100011110001001;
12'b110011111111: finv1 = 23'b00011010100001010101010;
12'b110100000000: finv1 = 23'b00011010011110111001011;
12'b110100000001: finv1 = 23'b00011010011100011101100;
12'b110100000010: finv1 = 23'b00011010011010000001110;
12'b110100000011: finv1 = 23'b00011010010111100110000;
12'b110100000100: finv1 = 23'b00011010010101001010010;
12'b110100000101: finv1 = 23'b00011010010010101110101;
12'b110100000110: finv1 = 23'b00011010010000010011000;
12'b110100000111: finv1 = 23'b00011010001101110111100;
12'b110100001000: finv1 = 23'b00011010001011011011111;
12'b110100001001: finv1 = 23'b00011010001001000000011;
12'b110100001010: finv1 = 23'b00011010000110100101000;
12'b110100001011: finv1 = 23'b00011010000100001001100;
12'b110100001100: finv1 = 23'b00011010000001101110001;
12'b110100001101: finv1 = 23'b00011001111111010010111;
12'b110100001110: finv1 = 23'b00011001111100110111100;
12'b110100001111: finv1 = 23'b00011001111010011100010;
12'b110100010000: finv1 = 23'b00011001111000000001001;
12'b110100010001: finv1 = 23'b00011001110101100110000;
12'b110100010010: finv1 = 23'b00011001110011001010111;
12'b110100010011: finv1 = 23'b00011001110000101111110;
12'b110100010100: finv1 = 23'b00011001101110010100110;
12'b110100010101: finv1 = 23'b00011001101011111001110;
12'b110100010110: finv1 = 23'b00011001101001011110110;
12'b110100010111: finv1 = 23'b00011001100111000011111;
12'b110100011000: finv1 = 23'b00011001100100101001000;
12'b110100011001: finv1 = 23'b00011001100010001110001;
12'b110100011010: finv1 = 23'b00011001011111110011011;
12'b110100011011: finv1 = 23'b00011001011101011000101;
12'b110100011100: finv1 = 23'b00011001011010111101111;
12'b110100011101: finv1 = 23'b00011001011000100011010;
12'b110100011110: finv1 = 23'b00011001010110001000101;
12'b110100011111: finv1 = 23'b00011001010011101110000;
12'b110100100000: finv1 = 23'b00011001010001010011100;
12'b110100100001: finv1 = 23'b00011001001110111001000;
12'b110100100010: finv1 = 23'b00011001001100011110100;
12'b110100100011: finv1 = 23'b00011001001010000100001;
12'b110100100100: finv1 = 23'b00011001000111101001110;
12'b110100100101: finv1 = 23'b00011001000101001111011;
12'b110100100110: finv1 = 23'b00011001000010110101001;
12'b110100100111: finv1 = 23'b00011001000000011010111;
12'b110100101000: finv1 = 23'b00011000111110000000101;
12'b110100101001: finv1 = 23'b00011000111011100110100;
12'b110100101010: finv1 = 23'b00011000111001001100011;
12'b110100101011: finv1 = 23'b00011000110110110010010;
12'b110100101100: finv1 = 23'b00011000110100011000010;
12'b110100101101: finv1 = 23'b00011000110001111110010;
12'b110100101110: finv1 = 23'b00011000101111100100010;
12'b110100101111: finv1 = 23'b00011000101101001010011;
12'b110100110000: finv1 = 23'b00011000101010110000100;
12'b110100110001: finv1 = 23'b00011000101000010110101;
12'b110100110010: finv1 = 23'b00011000100101111100111;
12'b110100110011: finv1 = 23'b00011000100011100011001;
12'b110100110100: finv1 = 23'b00011000100001001001011;
12'b110100110101: finv1 = 23'b00011000011110101111110;
12'b110100110110: finv1 = 23'b00011000011100010110001;
12'b110100110111: finv1 = 23'b00011000011001111100100;
12'b110100111000: finv1 = 23'b00011000010111100011000;
12'b110100111001: finv1 = 23'b00011000010101001001100;
12'b110100111010: finv1 = 23'b00011000010010110000000;
12'b110100111011: finv1 = 23'b00011000010000010110101;
12'b110100111100: finv1 = 23'b00011000001101111101010;
12'b110100111101: finv1 = 23'b00011000001011100011111;
12'b110100111110: finv1 = 23'b00011000001001001010100;
12'b110100111111: finv1 = 23'b00011000000110110001010;
12'b110101000000: finv1 = 23'b00011000000100011000001;
12'b110101000001: finv1 = 23'b00011000000001111110111;
12'b110101000010: finv1 = 23'b00010111111111100101110;
12'b110101000011: finv1 = 23'b00010111111101001100101;
12'b110101000100: finv1 = 23'b00010111111010110011101;
12'b110101000101: finv1 = 23'b00010111111000011010101;
12'b110101000110: finv1 = 23'b00010111110110000001101;
12'b110101000111: finv1 = 23'b00010111110011101000101;
12'b110101001000: finv1 = 23'b00010111110001001111110;
12'b110101001001: finv1 = 23'b00010111101110110110111;
12'b110101001010: finv1 = 23'b00010111101100011110001;
12'b110101001011: finv1 = 23'b00010111101010000101011;
12'b110101001100: finv1 = 23'b00010111100111101100101;
12'b110101001101: finv1 = 23'b00010111100101010011111;
12'b110101001110: finv1 = 23'b00010111100010111011010;
12'b110101001111: finv1 = 23'b00010111100000100010101;
12'b110101010000: finv1 = 23'b00010111011110001010001;
12'b110101010001: finv1 = 23'b00010111011011110001101;
12'b110101010010: finv1 = 23'b00010111011001011001001;
12'b110101010011: finv1 = 23'b00010111010111000000101;
12'b110101010100: finv1 = 23'b00010111010100101000010;
12'b110101010101: finv1 = 23'b00010111010010001111111;
12'b110101010110: finv1 = 23'b00010111001111110111100;
12'b110101010111: finv1 = 23'b00010111001101011111010;
12'b110101011000: finv1 = 23'b00010111001011000111000;
12'b110101011001: finv1 = 23'b00010111001000101110111;
12'b110101011010: finv1 = 23'b00010111000110010110101;
12'b110101011011: finv1 = 23'b00010111000011111110100;
12'b110101011100: finv1 = 23'b00010111000001100110100;
12'b110101011101: finv1 = 23'b00010110111111001110011;
12'b110101011110: finv1 = 23'b00010110111100110110011;
12'b110101011111: finv1 = 23'b00010110111010011110100;
12'b110101100000: finv1 = 23'b00010110111000000110100;
12'b110101100001: finv1 = 23'b00010110110101101110101;
12'b110101100010: finv1 = 23'b00010110110011010110111;
12'b110101100011: finv1 = 23'b00010110110000111111000;
12'b110101100100: finv1 = 23'b00010110101110100111010;
12'b110101100101: finv1 = 23'b00010110101100001111100;
12'b110101100110: finv1 = 23'b00010110101001110111111;
12'b110101100111: finv1 = 23'b00010110100111100000010;
12'b110101101000: finv1 = 23'b00010110100101001000101;
12'b110101101001: finv1 = 23'b00010110100010110001001;
12'b110101101010: finv1 = 23'b00010110100000011001101;
12'b110101101011: finv1 = 23'b00010110011110000010001;
12'b110101101100: finv1 = 23'b00010110011011101010101;
12'b110101101101: finv1 = 23'b00010110011001010011010;
12'b110101101110: finv1 = 23'b00010110010110111011111;
12'b110101101111: finv1 = 23'b00010110010100100100101;
12'b110101110000: finv1 = 23'b00010110010010001101011;
12'b110101110001: finv1 = 23'b00010110001111110110001;
12'b110101110010: finv1 = 23'b00010110001101011110111;
12'b110101110011: finv1 = 23'b00010110001011000111110;
12'b110101110100: finv1 = 23'b00010110001000110000101;
12'b110101110101: finv1 = 23'b00010110000110011001100;
12'b110101110110: finv1 = 23'b00010110000100000010100;
12'b110101110111: finv1 = 23'b00010110000001101011100;
12'b110101111000: finv1 = 23'b00010101111111010100101;
12'b110101111001: finv1 = 23'b00010101111100111101101;
12'b110101111010: finv1 = 23'b00010101111010100110110;
12'b110101111011: finv1 = 23'b00010101111000010000000;
12'b110101111100: finv1 = 23'b00010101110101111001001;
12'b110101111101: finv1 = 23'b00010101110011100010011;
12'b110101111110: finv1 = 23'b00010101110001001011101;
12'b110101111111: finv1 = 23'b00010101101110110101000;
12'b110110000000: finv1 = 23'b00010101101100011110011;
12'b110110000001: finv1 = 23'b00010101101010000111110;
12'b110110000010: finv1 = 23'b00010101100111110001010;
12'b110110000011: finv1 = 23'b00010101100101011010110;
12'b110110000100: finv1 = 23'b00010101100011000100010;
12'b110110000101: finv1 = 23'b00010101100000101101110;
12'b110110000110: finv1 = 23'b00010101011110010111011;
12'b110110000111: finv1 = 23'b00010101011100000001000;
12'b110110001000: finv1 = 23'b00010101011001101010110;
12'b110110001001: finv1 = 23'b00010101010111010100100;
12'b110110001010: finv1 = 23'b00010101010100111110010;
12'b110110001011: finv1 = 23'b00010101010010101000000;
12'b110110001100: finv1 = 23'b00010101010000010001111;
12'b110110001101: finv1 = 23'b00010101001101111011110;
12'b110110001110: finv1 = 23'b00010101001011100101101;
12'b110110001111: finv1 = 23'b00010101001001001111101;
12'b110110010000: finv1 = 23'b00010101000110111001101;
12'b110110010001: finv1 = 23'b00010101000100100011101;
12'b110110010010: finv1 = 23'b00010101000010001101110;
12'b110110010011: finv1 = 23'b00010100111111110111111;
12'b110110010100: finv1 = 23'b00010100111101100010000;
12'b110110010101: finv1 = 23'b00010100111011001100010;
12'b110110010110: finv1 = 23'b00010100111000110110100;
12'b110110010111: finv1 = 23'b00010100110110100000110;
12'b110110011000: finv1 = 23'b00010100110100001011001;
12'b110110011001: finv1 = 23'b00010100110001110101100;
12'b110110011010: finv1 = 23'b00010100101111011111111;
12'b110110011011: finv1 = 23'b00010100101101001010010;
12'b110110011100: finv1 = 23'b00010100101010110100110;
12'b110110011101: finv1 = 23'b00010100101000011111010;
12'b110110011110: finv1 = 23'b00010100100110001001111;
12'b110110011111: finv1 = 23'b00010100100011110100011;
12'b110110100000: finv1 = 23'b00010100100001011111000;
12'b110110100001: finv1 = 23'b00010100011111001001110;
12'b110110100010: finv1 = 23'b00010100011100110100100;
12'b110110100011: finv1 = 23'b00010100011010011111010;
12'b110110100100: finv1 = 23'b00010100011000001010000;
12'b110110100101: finv1 = 23'b00010100010101110100111;
12'b110110100110: finv1 = 23'b00010100010011011111110;
12'b110110100111: finv1 = 23'b00010100010001001010101;
12'b110110101000: finv1 = 23'b00010100001110110101100;
12'b110110101001: finv1 = 23'b00010100001100100000100;
12'b110110101010: finv1 = 23'b00010100001010001011101;
12'b110110101011: finv1 = 23'b00010100000111110110101;
12'b110110101100: finv1 = 23'b00010100000101100001110;
12'b110110101101: finv1 = 23'b00010100000011001100111;
12'b110110101110: finv1 = 23'b00010100000000111000001;
12'b110110101111: finv1 = 23'b00010011111110100011010;
12'b110110110000: finv1 = 23'b00010011111100001110100;
12'b110110110001: finv1 = 23'b00010011111001111001111;
12'b110110110010: finv1 = 23'b00010011110111100101010;
12'b110110110011: finv1 = 23'b00010011110101010000101;
12'b110110110100: finv1 = 23'b00010011110010111100000;
12'b110110110101: finv1 = 23'b00010011110000100111100;
12'b110110110110: finv1 = 23'b00010011101110010011000;
12'b110110110111: finv1 = 23'b00010011101011111110100;
12'b110110111000: finv1 = 23'b00010011101001101010000;
12'b110110111001: finv1 = 23'b00010011100111010101101;
12'b110110111010: finv1 = 23'b00010011100101000001011;
12'b110110111011: finv1 = 23'b00010011100010101101000;
12'b110110111100: finv1 = 23'b00010011100000011000110;
12'b110110111101: finv1 = 23'b00010011011110000100100;
12'b110110111110: finv1 = 23'b00010011011011110000011;
12'b110110111111: finv1 = 23'b00010011011001011100001;
12'b110111000000: finv1 = 23'b00010011010111001000001;
12'b110111000001: finv1 = 23'b00010011010100110100000;
12'b110111000010: finv1 = 23'b00010011010010100000000;
12'b110111000011: finv1 = 23'b00010011010000001100000;
12'b110111000100: finv1 = 23'b00010011001101111000000;
12'b110111000101: finv1 = 23'b00010011001011100100001;
12'b110111000110: finv1 = 23'b00010011001001010000010;
12'b110111000111: finv1 = 23'b00010011000110111100011;
12'b110111001000: finv1 = 23'b00010011000100101000100;
12'b110111001001: finv1 = 23'b00010011000010010100110;
12'b110111001010: finv1 = 23'b00010011000000000001001;
12'b110111001011: finv1 = 23'b00010010111101101101011;
12'b110111001100: finv1 = 23'b00010010111011011001110;
12'b110111001101: finv1 = 23'b00010010111001000110001;
12'b110111001110: finv1 = 23'b00010010110110110010101;
12'b110111001111: finv1 = 23'b00010010110100011111000;
12'b110111010000: finv1 = 23'b00010010110010001011100;
12'b110111010001: finv1 = 23'b00010010101111111000001;
12'b110111010010: finv1 = 23'b00010010101101100100101;
12'b110111010011: finv1 = 23'b00010010101011010001010;
12'b110111010100: finv1 = 23'b00010010101000111110000;
12'b110111010101: finv1 = 23'b00010010100110101010101;
12'b110111010110: finv1 = 23'b00010010100100010111011;
12'b110111010111: finv1 = 23'b00010010100010000100001;
12'b110111011000: finv1 = 23'b00010010011111110001000;
12'b110111011001: finv1 = 23'b00010010011101011101111;
12'b110111011010: finv1 = 23'b00010010011011001010110;
12'b110111011011: finv1 = 23'b00010010011000110111101;
12'b110111011100: finv1 = 23'b00010010010110100100101;
12'b110111011101: finv1 = 23'b00010010010100010001101;
12'b110111011110: finv1 = 23'b00010010010001111110110;
12'b110111011111: finv1 = 23'b00010010001111101011110;
12'b110111100000: finv1 = 23'b00010010001101011000111;
12'b110111100001: finv1 = 23'b00010010001011000110001;
12'b110111100010: finv1 = 23'b00010010001000110011010;
12'b110111100011: finv1 = 23'b00010010000110100000100;
12'b110111100100: finv1 = 23'b00010010000100001101110;
12'b110111100101: finv1 = 23'b00010010000001111011001;
12'b110111100110: finv1 = 23'b00010001111111101000100;
12'b110111100111: finv1 = 23'b00010001111101010101111;
12'b110111101000: finv1 = 23'b00010001111011000011010;
12'b110111101001: finv1 = 23'b00010001111000110000110;
12'b110111101010: finv1 = 23'b00010001110110011110010;
12'b110111101011: finv1 = 23'b00010001110100001011110;
12'b110111101100: finv1 = 23'b00010001110001111001011;
12'b110111101101: finv1 = 23'b00010001101111100111000;
12'b110111101110: finv1 = 23'b00010001101101010100101;
12'b110111101111: finv1 = 23'b00010001101011000010011;
12'b110111110000: finv1 = 23'b00010001101000110000001;
12'b110111110001: finv1 = 23'b00010001100110011101111;
12'b110111110010: finv1 = 23'b00010001100100001011110;
12'b110111110011: finv1 = 23'b00010001100001111001100;
12'b110111110100: finv1 = 23'b00010001011111100111011;
12'b110111110101: finv1 = 23'b00010001011101010101011;
12'b110111110110: finv1 = 23'b00010001011011000011011;
12'b110111110111: finv1 = 23'b00010001011000110001011;
12'b110111111000: finv1 = 23'b00010001010110011111011;
12'b110111111001: finv1 = 23'b00010001010100001101100;
12'b110111111010: finv1 = 23'b00010001010001111011101;
12'b110111111011: finv1 = 23'b00010001001111101001110;
12'b110111111100: finv1 = 23'b00010001001101010111111;
12'b110111111101: finv1 = 23'b00010001001011000110001;
12'b110111111110: finv1 = 23'b00010001001000110100011;
12'b110111111111: finv1 = 23'b00010001000110100010110;
12'b111000000000: finv1 = 23'b00010001000100010001001;
12'b111000000001: finv1 = 23'b00010001000001111111100;
12'b111000000010: finv1 = 23'b00010000111111101101111;
12'b111000000011: finv1 = 23'b00010000111101011100011;
12'b111000000100: finv1 = 23'b00010000111011001010111;
12'b111000000101: finv1 = 23'b00010000111000111001011;
12'b111000000110: finv1 = 23'b00010000110110100111111;
12'b111000000111: finv1 = 23'b00010000110100010110100;
12'b111000001000: finv1 = 23'b00010000110010000101010;
12'b111000001001: finv1 = 23'b00010000101111110011111;
12'b111000001010: finv1 = 23'b00010000101101100010101;
12'b111000001011: finv1 = 23'b00010000101011010001011;
12'b111000001100: finv1 = 23'b00010000101001000000001;
12'b111000001101: finv1 = 23'b00010000100110101111000;
12'b111000001110: finv1 = 23'b00010000100100011101111;
12'b111000001111: finv1 = 23'b00010000100010001100110;
12'b111000010000: finv1 = 23'b00010000011111111011110;
12'b111000010001: finv1 = 23'b00010000011101101010110;
12'b111000010010: finv1 = 23'b00010000011011011001110;
12'b111000010011: finv1 = 23'b00010000011001001000111;
12'b111000010100: finv1 = 23'b00010000010110110111111;
12'b111000010101: finv1 = 23'b00010000010100100111000;
12'b111000010110: finv1 = 23'b00010000010010010110010;
12'b111000010111: finv1 = 23'b00010000010000000101100;
12'b111000011000: finv1 = 23'b00010000001101110100110;
12'b111000011001: finv1 = 23'b00010000001011100100000;
12'b111000011010: finv1 = 23'b00010000001001010011011;
12'b111000011011: finv1 = 23'b00010000000111000010101;
12'b111000011100: finv1 = 23'b00010000000100110010001;
12'b111000011101: finv1 = 23'b00010000000010100001100;
12'b111000011110: finv1 = 23'b00010000000000010001000;
12'b111000011111: finv1 = 23'b00001111111110000000100;
12'b111000100000: finv1 = 23'b00001111111011110000001;
12'b111000100001: finv1 = 23'b00001111111001011111101;
12'b111000100010: finv1 = 23'b00001111110111001111010;
12'b111000100011: finv1 = 23'b00001111110100111111000;
12'b111000100100: finv1 = 23'b00001111110010101110101;
12'b111000100101: finv1 = 23'b00001111110000011110011;
12'b111000100110: finv1 = 23'b00001111101110001110001;
12'b111000100111: finv1 = 23'b00001111101011111110000;
12'b111000101000: finv1 = 23'b00001111101001101101111;
12'b111000101001: finv1 = 23'b00001111100111011101110;
12'b111000101010: finv1 = 23'b00001111100101001101101;
12'b111000101011: finv1 = 23'b00001111100010111101101;
12'b111000101100: finv1 = 23'b00001111100000101101101;
12'b111000101101: finv1 = 23'b00001111011110011101101;
12'b111000101110: finv1 = 23'b00001111011100001101110;
12'b111000101111: finv1 = 23'b00001111011001111101111;
12'b111000110000: finv1 = 23'b00001111010111101110000;
12'b111000110001: finv1 = 23'b00001111010101011110001;
12'b111000110010: finv1 = 23'b00001111010011001110011;
12'b111000110011: finv1 = 23'b00001111010000111110101;
12'b111000110100: finv1 = 23'b00001111001110101111000;
12'b111000110101: finv1 = 23'b00001111001100011111010;
12'b111000110110: finv1 = 23'b00001111001010001111101;
12'b111000110111: finv1 = 23'b00001111001000000000001;
12'b111000111000: finv1 = 23'b00001111000101110000100;
12'b111000111001: finv1 = 23'b00001111000011100001000;
12'b111000111010: finv1 = 23'b00001111000001010001100;
12'b111000111011: finv1 = 23'b00001110111111000010001;
12'b111000111100: finv1 = 23'b00001110111100110010101;
12'b111000111101: finv1 = 23'b00001110111010100011010;
12'b111000111110: finv1 = 23'b00001110111000010100000;
12'b111000111111: finv1 = 23'b00001110110110000100101;
12'b111001000000: finv1 = 23'b00001110110011110101011;
12'b111001000001: finv1 = 23'b00001110110001100110010;
12'b111001000010: finv1 = 23'b00001110101111010111000;
12'b111001000011: finv1 = 23'b00001110101101000111111;
12'b111001000100: finv1 = 23'b00001110101010111000110;
12'b111001000101: finv1 = 23'b00001110101000101001110;
12'b111001000110: finv1 = 23'b00001110100110011010101;
12'b111001000111: finv1 = 23'b00001110100100001011101;
12'b111001001000: finv1 = 23'b00001110100001111100110;
12'b111001001001: finv1 = 23'b00001110011111101101110;
12'b111001001010: finv1 = 23'b00001110011101011110111;
12'b111001001011: finv1 = 23'b00001110011011010000000;
12'b111001001100: finv1 = 23'b00001110011001000001010;
12'b111001001101: finv1 = 23'b00001110010110110010100;
12'b111001001110: finv1 = 23'b00001110010100100011110;
12'b111001001111: finv1 = 23'b00001110010010010101000;
12'b111001010000: finv1 = 23'b00001110010000000110011;
12'b111001010001: finv1 = 23'b00001110001101110111110;
12'b111001010010: finv1 = 23'b00001110001011101001001;
12'b111001010011: finv1 = 23'b00001110001001011010100;
12'b111001010100: finv1 = 23'b00001110000111001100000;
12'b111001010101: finv1 = 23'b00001110000100111101100;
12'b111001010110: finv1 = 23'b00001110000010101111001;
12'b111001010111: finv1 = 23'b00001110000000100000110;
12'b111001011000: finv1 = 23'b00001101111110010010011;
12'b111001011001: finv1 = 23'b00001101111100000100000;
12'b111001011010: finv1 = 23'b00001101111001110101110;
12'b111001011011: finv1 = 23'b00001101110111100111011;
12'b111001011100: finv1 = 23'b00001101110101011001010;
12'b111001011101: finv1 = 23'b00001101110011001011000;
12'b111001011110: finv1 = 23'b00001101110000111100111;
12'b111001011111: finv1 = 23'b00001101101110101110110;
12'b111001100000: finv1 = 23'b00001101101100100000101;
12'b111001100001: finv1 = 23'b00001101101010010010101;
12'b111001100010: finv1 = 23'b00001101101000000100101;
12'b111001100011: finv1 = 23'b00001101100101110110101;
12'b111001100100: finv1 = 23'b00001101100011101000110;
12'b111001100101: finv1 = 23'b00001101100001011010110;
12'b111001100110: finv1 = 23'b00001101011111001101000;
12'b111001100111: finv1 = 23'b00001101011100111111001;
12'b111001101000: finv1 = 23'b00001101011010110001011;
12'b111001101001: finv1 = 23'b00001101011000100011101;
12'b111001101010: finv1 = 23'b00001101010110010101111;
12'b111001101011: finv1 = 23'b00001101010100001000001;
12'b111001101100: finv1 = 23'b00001101010001111010100;
12'b111001101101: finv1 = 23'b00001101001111101100111;
12'b111001101110: finv1 = 23'b00001101001101011111011;
12'b111001101111: finv1 = 23'b00001101001011010001111;
12'b111001110000: finv1 = 23'b00001101001001000100011;
12'b111001110001: finv1 = 23'b00001101000110110110111;
12'b111001110010: finv1 = 23'b00001101000100101001100;
12'b111001110011: finv1 = 23'b00001101000010011100001;
12'b111001110100: finv1 = 23'b00001101000000001110110;
12'b111001110101: finv1 = 23'b00001100111110000001011;
12'b111001110110: finv1 = 23'b00001100111011110100001;
12'b111001110111: finv1 = 23'b00001100111001100110111;
12'b111001111000: finv1 = 23'b00001100110111011001101;
12'b111001111001: finv1 = 23'b00001100110101001100100;
12'b111001111010: finv1 = 23'b00001100110010111111011;
12'b111001111011: finv1 = 23'b00001100110000110010010;
12'b111001111100: finv1 = 23'b00001100101110100101010;
12'b111001111101: finv1 = 23'b00001100101100011000001;
12'b111001111110: finv1 = 23'b00001100101010001011001;
12'b111001111111: finv1 = 23'b00001100100111111110010;
12'b111010000000: finv1 = 23'b00001100100101110001010;
12'b111010000001: finv1 = 23'b00001100100011100100011;
12'b111010000010: finv1 = 23'b00001100100001010111101;
12'b111010000011: finv1 = 23'b00001100011111001010110;
12'b111010000100: finv1 = 23'b00001100011100111110000;
12'b111010000101: finv1 = 23'b00001100011010110001010;
12'b111010000110: finv1 = 23'b00001100011000100100100;
12'b111010000111: finv1 = 23'b00001100010110010111111;
12'b111010001000: finv1 = 23'b00001100010100001011010;
12'b111010001001: finv1 = 23'b00001100010001111110101;
12'b111010001010: finv1 = 23'b00001100001111110010001;
12'b111010001011: finv1 = 23'b00001100001101100101101;
12'b111010001100: finv1 = 23'b00001100001011011001001;
12'b111010001101: finv1 = 23'b00001100001001001100101;
12'b111010001110: finv1 = 23'b00001100000111000000010;
12'b111010001111: finv1 = 23'b00001100000100110011111;
12'b111010010000: finv1 = 23'b00001100000010100111100;
12'b111010010001: finv1 = 23'b00001100000000011011010;
12'b111010010010: finv1 = 23'b00001011111110001111000;
12'b111010010011: finv1 = 23'b00001011111100000010110;
12'b111010010100: finv1 = 23'b00001011111001110110100;
12'b111010010101: finv1 = 23'b00001011110111101010011;
12'b111010010110: finv1 = 23'b00001011110101011110010;
12'b111010010111: finv1 = 23'b00001011110011010010001;
12'b111010011000: finv1 = 23'b00001011110001000110001;
12'b111010011001: finv1 = 23'b00001011101110111010000;
12'b111010011010: finv1 = 23'b00001011101100101110001;
12'b111010011011: finv1 = 23'b00001011101010100010001;
12'b111010011100: finv1 = 23'b00001011101000010110010;
12'b111010011101: finv1 = 23'b00001011100110001010011;
12'b111010011110: finv1 = 23'b00001011100011111110100;
12'b111010011111: finv1 = 23'b00001011100001110010110;
12'b111010100000: finv1 = 23'b00001011011111100110111;
12'b111010100001: finv1 = 23'b00001011011101011011010;
12'b111010100010: finv1 = 23'b00001011011011001111100;
12'b111010100011: finv1 = 23'b00001011011001000011111;
12'b111010100100: finv1 = 23'b00001011010110111000010;
12'b111010100101: finv1 = 23'b00001011010100101100101;
12'b111010100110: finv1 = 23'b00001011010010100001000;
12'b111010100111: finv1 = 23'b00001011010000010101100;
12'b111010101000: finv1 = 23'b00001011001110001010000;
12'b111010101001: finv1 = 23'b00001011001011111110101;
12'b111010101010: finv1 = 23'b00001011001001110011001;
12'b111010101011: finv1 = 23'b00001011000111100111110;
12'b111010101100: finv1 = 23'b00001011000101011100100;
12'b111010101101: finv1 = 23'b00001011000011010001001;
12'b111010101110: finv1 = 23'b00001011000001000101111;
12'b111010101111: finv1 = 23'b00001010111110111010101;
12'b111010110000: finv1 = 23'b00001010111100101111100;
12'b111010110001: finv1 = 23'b00001010111010100100010;
12'b111010110010: finv1 = 23'b00001010111000011001001;
12'b111010110011: finv1 = 23'b00001010110110001110000;
12'b111010110100: finv1 = 23'b00001010110100000011000;
12'b111010110101: finv1 = 23'b00001010110001111000000;
12'b111010110110: finv1 = 23'b00001010101111101101000;
12'b111010110111: finv1 = 23'b00001010101101100010000;
12'b111010111000: finv1 = 23'b00001010101011010111001;
12'b111010111001: finv1 = 23'b00001010101001001100010;
12'b111010111010: finv1 = 23'b00001010100111000001011;
12'b111010111011: finv1 = 23'b00001010100100110110101;
12'b111010111100: finv1 = 23'b00001010100010101011110;
12'b111010111101: finv1 = 23'b00001010100000100001000;
12'b111010111110: finv1 = 23'b00001010011110010110011;
12'b111010111111: finv1 = 23'b00001010011100001011101;
12'b111011000000: finv1 = 23'b00001010011010000001000;
12'b111011000001: finv1 = 23'b00001010010111110110100;
12'b111011000010: finv1 = 23'b00001010010101101011111;
12'b111011000011: finv1 = 23'b00001010010011100001011;
12'b111011000100: finv1 = 23'b00001010010001010110111;
12'b111011000101: finv1 = 23'b00001010001111001100011;
12'b111011000110: finv1 = 23'b00001010001101000010000;
12'b111011000111: finv1 = 23'b00001010001010110111101;
12'b111011001000: finv1 = 23'b00001010001000101101010;
12'b111011001001: finv1 = 23'b00001010000110100010111;
12'b111011001010: finv1 = 23'b00001010000100011000101;
12'b111011001011: finv1 = 23'b00001010000010001110011;
12'b111011001100: finv1 = 23'b00001010000000000100001;
12'b111011001101: finv1 = 23'b00001001111101111010000;
12'b111011001110: finv1 = 23'b00001001111011101111111;
12'b111011001111: finv1 = 23'b00001001111001100101110;
12'b111011010000: finv1 = 23'b00001001110111011011101;
12'b111011010001: finv1 = 23'b00001001110101010001101;
12'b111011010010: finv1 = 23'b00001001110011000111101;
12'b111011010011: finv1 = 23'b00001001110000111101101;
12'b111011010100: finv1 = 23'b00001001101110110011110;
12'b111011010101: finv1 = 23'b00001001101100101001110;
12'b111011010110: finv1 = 23'b00001001101010100000000;
12'b111011010111: finv1 = 23'b00001001101000010110001;
12'b111011011000: finv1 = 23'b00001001100110001100011;
12'b111011011001: finv1 = 23'b00001001100100000010100;
12'b111011011010: finv1 = 23'b00001001100001111000111;
12'b111011011011: finv1 = 23'b00001001011111101111001;
12'b111011011100: finv1 = 23'b00001001011101100101100;
12'b111011011101: finv1 = 23'b00001001011011011011111;
12'b111011011110: finv1 = 23'b00001001011001010010010;
12'b111011011111: finv1 = 23'b00001001010111001000110;
12'b111011100000: finv1 = 23'b00001001010100111111010;
12'b111011100001: finv1 = 23'b00001001010010110101110;
12'b111011100010: finv1 = 23'b00001001010000101100010;
12'b111011100011: finv1 = 23'b00001001001110100010111;
12'b111011100100: finv1 = 23'b00001001001100011001100;
12'b111011100101: finv1 = 23'b00001001001010010000001;
12'b111011100110: finv1 = 23'b00001001001000000110111;
12'b111011100111: finv1 = 23'b00001001000101111101101;
12'b111011101000: finv1 = 23'b00001001000011110100011;
12'b111011101001: finv1 = 23'b00001001000001101011001;
12'b111011101010: finv1 = 23'b00001000111111100010000;
12'b111011101011: finv1 = 23'b00001000111101011000111;
12'b111011101100: finv1 = 23'b00001000111011001111110;
12'b111011101101: finv1 = 23'b00001000111001000110101;
12'b111011101110: finv1 = 23'b00001000110110111101101;
12'b111011101111: finv1 = 23'b00001000110100110100101;
12'b111011110000: finv1 = 23'b00001000110010101011110;
12'b111011110001: finv1 = 23'b00001000110000100010110;
12'b111011110010: finv1 = 23'b00001000101110011001111;
12'b111011110011: finv1 = 23'b00001000101100010001000;
12'b111011110100: finv1 = 23'b00001000101010001000010;
12'b111011110101: finv1 = 23'b00001000100111111111011;
12'b111011110110: finv1 = 23'b00001000100101110110101;
12'b111011110111: finv1 = 23'b00001000100011101110000;
12'b111011111000: finv1 = 23'b00001000100001100101010;
12'b111011111001: finv1 = 23'b00001000011111011100101;
12'b111011111010: finv1 = 23'b00001000011101010100000;
12'b111011111011: finv1 = 23'b00001000011011001011011;
12'b111011111100: finv1 = 23'b00001000011001000010111;
12'b111011111101: finv1 = 23'b00001000010110111010011;
12'b111011111110: finv1 = 23'b00001000010100110001111;
12'b111011111111: finv1 = 23'b00001000010010101001100;
12'b111100000000: finv1 = 23'b00001000010000100001000;
12'b111100000001: finv1 = 23'b00001000001110011000101;
12'b111100000010: finv1 = 23'b00001000001100010000011;
12'b111100000011: finv1 = 23'b00001000001010001000000;
12'b111100000100: finv1 = 23'b00001000000111111111110;
12'b111100000101: finv1 = 23'b00001000000101110111100;
12'b111100000110: finv1 = 23'b00001000000011101111010;
12'b111100000111: finv1 = 23'b00001000000001100111001;
12'b111100001000: finv1 = 23'b00000111111111011111000;
12'b111100001001: finv1 = 23'b00000111111101010110111;
12'b111100001010: finv1 = 23'b00000111111011001110111;
12'b111100001011: finv1 = 23'b00000111111001000110110;
12'b111100001100: finv1 = 23'b00000111110110111110110;
12'b111100001101: finv1 = 23'b00000111110100110110111;
12'b111100001110: finv1 = 23'b00000111110010101110111;
12'b111100001111: finv1 = 23'b00000111110000100111000;
12'b111100010000: finv1 = 23'b00000111101110011111001;
12'b111100010001: finv1 = 23'b00000111101100010111011;
12'b111100010010: finv1 = 23'b00000111101010001111100;
12'b111100010011: finv1 = 23'b00000111101000000111110;
12'b111100010100: finv1 = 23'b00000111100110000000001;
12'b111100010101: finv1 = 23'b00000111100011111000011;
12'b111100010110: finv1 = 23'b00000111100001110000110;
12'b111100010111: finv1 = 23'b00000111011111101001001;
12'b111100011000: finv1 = 23'b00000111011101100001100;
12'b111100011001: finv1 = 23'b00000111011011011010000;
12'b111100011010: finv1 = 23'b00000111011001010010100;
12'b111100011011: finv1 = 23'b00000111010111001011000;
12'b111100011100: finv1 = 23'b00000111010101000011100;
12'b111100011101: finv1 = 23'b00000111010010111100001;
12'b111100011110: finv1 = 23'b00000111010000110100110;
12'b111100011111: finv1 = 23'b00000111001110101101011;
12'b111100100000: finv1 = 23'b00000111001100100110000;
12'b111100100001: finv1 = 23'b00000111001010011110110;
12'b111100100010: finv1 = 23'b00000111001000010111100;
12'b111100100011: finv1 = 23'b00000111000110010000010;
12'b111100100100: finv1 = 23'b00000111000100001001001;
12'b111100100101: finv1 = 23'b00000111000010000010000;
12'b111100100110: finv1 = 23'b00000110111111111010111;
12'b111100100111: finv1 = 23'b00000110111101110011110;
12'b111100101000: finv1 = 23'b00000110111011101100110;
12'b111100101001: finv1 = 23'b00000110111001100101110;
12'b111100101010: finv1 = 23'b00000110110111011110110;
12'b111100101011: finv1 = 23'b00000110110101010111111;
12'b111100101100: finv1 = 23'b00000110110011010000111;
12'b111100101101: finv1 = 23'b00000110110001001010000;
12'b111100101110: finv1 = 23'b00000110101111000011010;
12'b111100101111: finv1 = 23'b00000110101100111100011;
12'b111100110000: finv1 = 23'b00000110101010110101101;
12'b111100110001: finv1 = 23'b00000110101000101110111;
12'b111100110010: finv1 = 23'b00000110100110101000001;
12'b111100110011: finv1 = 23'b00000110100100100001100;
12'b111100110100: finv1 = 23'b00000110100010011010111;
12'b111100110101: finv1 = 23'b00000110100000010100010;
12'b111100110110: finv1 = 23'b00000110011110001101101;
12'b111100110111: finv1 = 23'b00000110011100000111001;
12'b111100111000: finv1 = 23'b00000110011010000000101;
12'b111100111001: finv1 = 23'b00000110010111111010001;
12'b111100111010: finv1 = 23'b00000110010101110011110;
12'b111100111011: finv1 = 23'b00000110010011101101011;
12'b111100111100: finv1 = 23'b00000110010001100111000;
12'b111100111101: finv1 = 23'b00000110001111100000101;
12'b111100111110: finv1 = 23'b00000110001101011010011;
12'b111100111111: finv1 = 23'b00000110001011010100000;
12'b111101000000: finv1 = 23'b00000110001001001101111;
12'b111101000001: finv1 = 23'b00000110000111000111101;
12'b111101000010: finv1 = 23'b00000110000101000001100;
12'b111101000011: finv1 = 23'b00000110000010111011011;
12'b111101000100: finv1 = 23'b00000110000000110101010;
12'b111101000101: finv1 = 23'b00000101111110101111001;
12'b111101000110: finv1 = 23'b00000101111100101001001;
12'b111101000111: finv1 = 23'b00000101111010100011001;
12'b111101001000: finv1 = 23'b00000101111000011101001;
12'b111101001001: finv1 = 23'b00000101110110010111010;
12'b111101001010: finv1 = 23'b00000101110100010001011;
12'b111101001011: finv1 = 23'b00000101110010001011100;
12'b111101001100: finv1 = 23'b00000101110000000101101;
12'b111101001101: finv1 = 23'b00000101101101111111111;
12'b111101001110: finv1 = 23'b00000101101011111010000;
12'b111101001111: finv1 = 23'b00000101101001110100011;
12'b111101010000: finv1 = 23'b00000101100111101110101;
12'b111101010001: finv1 = 23'b00000101100101101001000;
12'b111101010010: finv1 = 23'b00000101100011100011011;
12'b111101010011: finv1 = 23'b00000101100001011101110;
12'b111101010100: finv1 = 23'b00000101011111011000001;
12'b111101010101: finv1 = 23'b00000101011101010010101;
12'b111101010110: finv1 = 23'b00000101011011001101001;
12'b111101010111: finv1 = 23'b00000101011001000111101;
12'b111101011000: finv1 = 23'b00000101010111000010010;
12'b111101011001: finv1 = 23'b00000101010100111100111;
12'b111101011010: finv1 = 23'b00000101010010110111100;
12'b111101011011: finv1 = 23'b00000101010000110010001;
12'b111101011100: finv1 = 23'b00000101001110101100111;
12'b111101011101: finv1 = 23'b00000101001100100111101;
12'b111101011110: finv1 = 23'b00000101001010100010011;
12'b111101011111: finv1 = 23'b00000101001000011101001;
12'b111101100000: finv1 = 23'b00000101000110011000000;
12'b111101100001: finv1 = 23'b00000101000100010010111;
12'b111101100010: finv1 = 23'b00000101000010001101110;
12'b111101100011: finv1 = 23'b00000101000000001000101;
12'b111101100100: finv1 = 23'b00000100111110000011101;
12'b111101100101: finv1 = 23'b00000100111011111110101;
12'b111101100110: finv1 = 23'b00000100111001111001101;
12'b111101100111: finv1 = 23'b00000100110111110100110;
12'b111101101000: finv1 = 23'b00000100110101101111111;
12'b111101101001: finv1 = 23'b00000100110011101011000;
12'b111101101010: finv1 = 23'b00000100110001100110001;
12'b111101101011: finv1 = 23'b00000100101111100001011;
12'b111101101100: finv1 = 23'b00000100101101011100100;
12'b111101101101: finv1 = 23'b00000100101011010111110;
12'b111101101110: finv1 = 23'b00000100101001010011001;
12'b111101101111: finv1 = 23'b00000100100111001110011;
12'b111101110000: finv1 = 23'b00000100100101001001110;
12'b111101110001: finv1 = 23'b00000100100011000101010;
12'b111101110010: finv1 = 23'b00000100100001000000101;
12'b111101110011: finv1 = 23'b00000100011110111100001;
12'b111101110100: finv1 = 23'b00000100011100110111101;
12'b111101110101: finv1 = 23'b00000100011010110011001;
12'b111101110110: finv1 = 23'b00000100011000101110101;
12'b111101110111: finv1 = 23'b00000100010110101010010;
12'b111101111000: finv1 = 23'b00000100010100100101111;
12'b111101111001: finv1 = 23'b00000100010010100001100;
12'b111101111010: finv1 = 23'b00000100010000011101010;
12'b111101111011: finv1 = 23'b00000100001110011001000;
12'b111101111100: finv1 = 23'b00000100001100010100110;
12'b111101111101: finv1 = 23'b00000100001010010000100;
12'b111101111110: finv1 = 23'b00000100001000001100011;
12'b111101111111: finv1 = 23'b00000100000110001000001;
12'b111110000000: finv1 = 23'b00000100000100000100001;
12'b111110000001: finv1 = 23'b00000100000010000000000;
12'b111110000010: finv1 = 23'b00000011111111111100000;
12'b111110000011: finv1 = 23'b00000011111101110111111;
12'b111110000100: finv1 = 23'b00000011111011110100000;
12'b111110000101: finv1 = 23'b00000011111001110000000;
12'b111110000110: finv1 = 23'b00000011110111101100001;
12'b111110000111: finv1 = 23'b00000011110101101000010;
12'b111110001000: finv1 = 23'b00000011110011100100011;
12'b111110001001: finv1 = 23'b00000011110001100000100;
12'b111110001010: finv1 = 23'b00000011101111011100110;
12'b111110001011: finv1 = 23'b00000011101101011001000;
12'b111110001100: finv1 = 23'b00000011101011010101010;
12'b111110001101: finv1 = 23'b00000011101001010001101;
12'b111110001110: finv1 = 23'b00000011100111001101111;
12'b111110001111: finv1 = 23'b00000011100101001010010;
12'b111110010000: finv1 = 23'b00000011100011000110110;
12'b111110010001: finv1 = 23'b00000011100001000011001;
12'b111110010010: finv1 = 23'b00000011011110111111101;
12'b111110010011: finv1 = 23'b00000011011100111100001;
12'b111110010100: finv1 = 23'b00000011011010111000101;
12'b111110010101: finv1 = 23'b00000011011000110101010;
12'b111110010110: finv1 = 23'b00000011010110110001111;
12'b111110010111: finv1 = 23'b00000011010100101110100;
12'b111110011000: finv1 = 23'b00000011010010101011001;
12'b111110011001: finv1 = 23'b00000011010000100111111;
12'b111110011010: finv1 = 23'b00000011001110100100101;
12'b111110011011: finv1 = 23'b00000011001100100001011;
12'b111110011100: finv1 = 23'b00000011001010011110001;
12'b111110011101: finv1 = 23'b00000011001000011011000;
12'b111110011110: finv1 = 23'b00000011000110010111111;
12'b111110011111: finv1 = 23'b00000011000100010100110;
12'b111110100000: finv1 = 23'b00000011000010010001110;
12'b111110100001: finv1 = 23'b00000011000000001110101;
12'b111110100010: finv1 = 23'b00000010111110001011101;
12'b111110100011: finv1 = 23'b00000010111100001000110;
12'b111110100100: finv1 = 23'b00000010111010000101110;
12'b111110100101: finv1 = 23'b00000010111000000010111;
12'b111110100110: finv1 = 23'b00000010110110000000000;
12'b111110100111: finv1 = 23'b00000010110011111101001;
12'b111110101000: finv1 = 23'b00000010110001111010011;
12'b111110101001: finv1 = 23'b00000010101111110111100;
12'b111110101010: finv1 = 23'b00000010101101110100110;
12'b111110101011: finv1 = 23'b00000010101011110010001;
12'b111110101100: finv1 = 23'b00000010101001101111011;
12'b111110101101: finv1 = 23'b00000010100111101100110;
12'b111110101110: finv1 = 23'b00000010100101101010001;
12'b111110101111: finv1 = 23'b00000010100011100111100;
12'b111110110000: finv1 = 23'b00000010100001100101000;
12'b111110110001: finv1 = 23'b00000010011111100010100;
12'b111110110010: finv1 = 23'b00000010011101100000000;
12'b111110110011: finv1 = 23'b00000010011011011101100;
12'b111110110100: finv1 = 23'b00000010011001011011001;
12'b111110110101: finv1 = 23'b00000010010111011000110;
12'b111110110110: finv1 = 23'b00000010010101010110011;
12'b111110110111: finv1 = 23'b00000010010011010100000;
12'b111110111000: finv1 = 23'b00000010010001010001110;
12'b111110111001: finv1 = 23'b00000010001111001111100;
12'b111110111010: finv1 = 23'b00000010001101001101010;
12'b111110111011: finv1 = 23'b00000010001011001011000;
12'b111110111100: finv1 = 23'b00000010001001001000111;
12'b111110111101: finv1 = 23'b00000010000111000110110;
12'b111110111110: finv1 = 23'b00000010000101000100101;
12'b111110111111: finv1 = 23'b00000010000011000010100;
12'b111111000000: finv1 = 23'b00000010000001000000100;
12'b111111000001: finv1 = 23'b00000001111110111110100;
12'b111111000010: finv1 = 23'b00000001111100111100100;
12'b111111000011: finv1 = 23'b00000001111010111010101;
12'b111111000100: finv1 = 23'b00000001111000111000101;
12'b111111000101: finv1 = 23'b00000001110110110110110;
12'b111111000110: finv1 = 23'b00000001110100110100111;
12'b111111000111: finv1 = 23'b00000001110010110011001;
12'b111111001000: finv1 = 23'b00000001110000110001011;
12'b111111001001: finv1 = 23'b00000001101110101111101;
12'b111111001010: finv1 = 23'b00000001101100101101111;
12'b111111001011: finv1 = 23'b00000001101010101100001;
12'b111111001100: finv1 = 23'b00000001101000101010100;
12'b111111001101: finv1 = 23'b00000001100110101000111;
12'b111111001110: finv1 = 23'b00000001100100100111010;
12'b111111001111: finv1 = 23'b00000001100010100101110;
12'b111111010000: finv1 = 23'b00000001100000100100010;
12'b111111010001: finv1 = 23'b00000001011110100010110;
12'b111111010010: finv1 = 23'b00000001011100100001010;
12'b111111010011: finv1 = 23'b00000001011010011111111;
12'b111111010100: finv1 = 23'b00000001011000011110011;
12'b111111010101: finv1 = 23'b00000001010110011101000;
12'b111111010110: finv1 = 23'b00000001010100011011110;
12'b111111010111: finv1 = 23'b00000001010010011010011;
12'b111111011000: finv1 = 23'b00000001010000011001001;
12'b111111011001: finv1 = 23'b00000001001110010111111;
12'b111111011010: finv1 = 23'b00000001001100010110101;
12'b111111011011: finv1 = 23'b00000001001010010101100;
12'b111111011100: finv1 = 23'b00000001001000010100011;
12'b111111011101: finv1 = 23'b00000001000110010011010;
12'b111111011110: finv1 = 23'b00000001000100010010001;
12'b111111011111: finv1 = 23'b00000001000010010001001;
12'b111111100000: finv1 = 23'b00000001000000010000001;
12'b111111100001: finv1 = 23'b00000000111110001111001;
12'b111111100010: finv1 = 23'b00000000111100001110001;
12'b111111100011: finv1 = 23'b00000000111010001101001;
12'b111111100100: finv1 = 23'b00000000111000001100010;
12'b111111100101: finv1 = 23'b00000000110110001011011;
12'b111111100110: finv1 = 23'b00000000110100001010101;
12'b111111100111: finv1 = 23'b00000000110010001001110;
12'b111111101000: finv1 = 23'b00000000110000001001000;
12'b111111101001: finv1 = 23'b00000000101110001000010;
12'b111111101010: finv1 = 23'b00000000101100000111101;
12'b111111101011: finv1 = 23'b00000000101010000110111;
12'b111111101100: finv1 = 23'b00000000101000000110010;
12'b111111101101: finv1 = 23'b00000000100110000101101;
12'b111111101110: finv1 = 23'b00000000100100000101001;
12'b111111101111: finv1 = 23'b00000000100010000100100;
12'b111111110000: finv1 = 23'b00000000100000000100000;
12'b111111110001: finv1 = 23'b00000000011110000011100;
12'b111111110010: finv1 = 23'b00000000011100000011001;
12'b111111110011: finv1 = 23'b00000000011010000010101;
12'b111111110100: finv1 = 23'b00000000011000000010010;
12'b111111110101: finv1 = 23'b00000000010110000001111;
12'b111111110110: finv1 = 23'b00000000010100000001101;
12'b111111110111: finv1 = 23'b00000000010010000001010;
12'b111111111000: finv1 = 23'b00000000010000000001000;
12'b111111111001: finv1 = 23'b00000000001110000000110;
12'b111111111010: finv1 = 23'b00000000001100000000101;
12'b111111111011: finv1 = 23'b00000000001010000000011;
12'b111111111100: finv1 = 23'b00000000001000000000010;
12'b111111111101: finv1 = 23'b00000000000110000000001;
12'b111111111110: finv1 = 23'b00000000000100000000001;
12'b111111111111: finv1 = 23'b00000000000010000000000;

     endcase
    end
  endfunction

  function [22:0] finv2 (
    input [11:0] m_input2 );
    begin
      case(m_input2)

12'b000000000000: finv2 = 23'b00000000000000000000000;
12'b000000000001: finv2 = 23'b11111111110000000000011;
12'b000000000010: finv2 = 23'b11111111100000000001100;
12'b000000000011: finv2 = 23'b11111111010000000011011;
12'b000000000100: finv2 = 23'b11111111000000000110000;
12'b000000000101: finv2 = 23'b11111110110000001001011;
12'b000000000110: finv2 = 23'b11111110100000001101100;
12'b000000000111: finv2 = 23'b11111110010000010010011;
12'b000000001000: finv2 = 23'b11111110000000011000000;
12'b000000001001: finv2 = 23'b11111101110000011110010;
12'b000000001010: finv2 = 23'b11111101100000100101011;
12'b000000001011: finv2 = 23'b11111101010000101101010;
12'b000000001100: finv2 = 23'b11111101000000110101110;
12'b000000001101: finv2 = 23'b11111100110000111111001;
12'b000000001110: finv2 = 23'b11111100100001001001001;
12'b000000001111: finv2 = 23'b11111100010001010100000;
12'b000000010000: finv2 = 23'b11111100000001011111100;
12'b000000010001: finv2 = 23'b11111011110001101011110;
12'b000000010010: finv2 = 23'b11111011100001111000110;
12'b000000010011: finv2 = 23'b11111011010010000110100;
12'b000000010100: finv2 = 23'b11111011000010010101000;
12'b000000010101: finv2 = 23'b11111010110010100100010;
12'b000000010110: finv2 = 23'b11111010100010110100010;
12'b000000010111: finv2 = 23'b11111010010011000100111;
12'b000000011000: finv2 = 23'b11111010000011010110011;
12'b000000011001: finv2 = 23'b11111001110011101000100;
12'b000000011010: finv2 = 23'b11111001100011111011011;
12'b000000011011: finv2 = 23'b11111001010100001111000;
12'b000000011100: finv2 = 23'b11111001000100100011011;
12'b000000011101: finv2 = 23'b11111000110100111000011;
12'b000000011110: finv2 = 23'b11111000100101001110010;
12'b000000011111: finv2 = 23'b11111000010101100100110;
12'b000000100000: finv2 = 23'b11111000000101111100000;
12'b000000100001: finv2 = 23'b11110111110110010100000;
12'b000000100010: finv2 = 23'b11110111100110101100110;
12'b000000100011: finv2 = 23'b11110111010111000110010;
12'b000000100100: finv2 = 23'b11110111000111100000011;
12'b000000100101: finv2 = 23'b11110110110111111011010;
12'b000000100110: finv2 = 23'b11110110101000010110111;
12'b000000100111: finv2 = 23'b11110110011000110011010;
12'b000000101000: finv2 = 23'b11110110001001010000010;
12'b000000101001: finv2 = 23'b11110101111001101110001;
12'b000000101010: finv2 = 23'b11110101101010001100101;
12'b000000101011: finv2 = 23'b11110101011010101011110;
12'b000000101100: finv2 = 23'b11110101001011001011110;
12'b000000101101: finv2 = 23'b11110100111011101100011;
12'b000000101110: finv2 = 23'b11110100101100001101110;
12'b000000101111: finv2 = 23'b11110100011100101111111;
12'b000000110000: finv2 = 23'b11110100001101010010110;
12'b000000110001: finv2 = 23'b11110011111101110110010;
12'b000000110010: finv2 = 23'b11110011101110011010100;
12'b000000110011: finv2 = 23'b11110011011110111111011;
12'b000000110100: finv2 = 23'b11110011001111100101001;
12'b000000110101: finv2 = 23'b11110011000000001011100;
12'b000000110110: finv2 = 23'b11110010110000110010101;
12'b000000110111: finv2 = 23'b11110010100001011010011;
12'b000000111000: finv2 = 23'b11110010010010000010111;
12'b000000111001: finv2 = 23'b11110010000010101100001;
12'b000000111010: finv2 = 23'b11110001110011010110001;
12'b000000111011: finv2 = 23'b11110001100100000000110;
12'b000000111100: finv2 = 23'b11110001010100101100001;
12'b000000111101: finv2 = 23'b11110001000101011000001;
12'b000000111110: finv2 = 23'b11110000110110000101000;
12'b000000111111: finv2 = 23'b11110000100110110010011;
12'b000001000000: finv2 = 23'b11110000010111100000101;
12'b000001000001: finv2 = 23'b11110000001000001111100;
12'b000001000010: finv2 = 23'b11101111111000111111001;
12'b000001000011: finv2 = 23'b11101111101001101111011;
12'b000001000100: finv2 = 23'b11101111011010100000011;
12'b000001000101: finv2 = 23'b11101111001011010010001;
12'b000001000110: finv2 = 23'b11101110111100000100100;
12'b000001000111: finv2 = 23'b11101110101100110111101;
12'b000001001000: finv2 = 23'b11101110011101101011011;
12'b000001001001: finv2 = 23'b11101110001110011111111;
12'b000001001010: finv2 = 23'b11101101111111010101001;
12'b000001001011: finv2 = 23'b11101101110000001011000;
12'b000001001100: finv2 = 23'b11101101100001000001101;
12'b000001001101: finv2 = 23'b11101101010001111000111;
12'b000001001110: finv2 = 23'b11101101000010110000111;
12'b000001001111: finv2 = 23'b11101100110011101001101;
12'b000001010000: finv2 = 23'b11101100100100100011000;
12'b000001010001: finv2 = 23'b11101100010101011101001;
12'b000001010010: finv2 = 23'b11101100000110010111111;
12'b000001010011: finv2 = 23'b11101011110111010011010;
12'b000001010100: finv2 = 23'b11101011101000001111100;
12'b000001010101: finv2 = 23'b11101011011001001100010;
12'b000001010110: finv2 = 23'b11101011001010001001111;
12'b000001010111: finv2 = 23'b11101010111011001000001;
12'b000001011000: finv2 = 23'b11101010101100000111000;
12'b000001011001: finv2 = 23'b11101010011101000110101;
12'b000001011010: finv2 = 23'b11101010001110000110111;
12'b000001011011: finv2 = 23'b11101001111111000111111;
12'b000001011100: finv2 = 23'b11101001110000001001100;
12'b000001011101: finv2 = 23'b11101001100001001011111;
12'b000001011110: finv2 = 23'b11101001010010001111000;
12'b000001011111: finv2 = 23'b11101001000011010010101;
12'b000001100000: finv2 = 23'b11101000110100010111001;
12'b000001100001: finv2 = 23'b11101000100101011100001;
12'b000001100010: finv2 = 23'b11101000010110100010000;
12'b000001100011: finv2 = 23'b11101000000111101000011;
12'b000001100100: finv2 = 23'b11100111111000101111100;
12'b000001100101: finv2 = 23'b11100111101001110111011;
12'b000001100110: finv2 = 23'b11100111011010111111111;
12'b000001100111: finv2 = 23'b11100111001100001001000;
12'b000001101000: finv2 = 23'b11100110111101010010111;
12'b000001101001: finv2 = 23'b11100110101110011101100;
12'b000001101010: finv2 = 23'b11100110011111101000101;
12'b000001101011: finv2 = 23'b11100110010000110100101;
12'b000001101100: finv2 = 23'b11100110000010000001001;
12'b000001101101: finv2 = 23'b11100101110011001110011;
12'b000001101110: finv2 = 23'b11100101100100011100010;
12'b000001101111: finv2 = 23'b11100101010101101010111;
12'b000001110000: finv2 = 23'b11100101000110111010001;
12'b000001110001: finv2 = 23'b11100100111000001010001;
12'b000001110010: finv2 = 23'b11100100101001011010110;
12'b000001110011: finv2 = 23'b11100100011010101100000;
12'b000001110100: finv2 = 23'b11100100001011111110000;
12'b000001110101: finv2 = 23'b11100011111101010000101;
12'b000001110110: finv2 = 23'b11100011101110100011111;
12'b000001110111: finv2 = 23'b11100011011111110111111;
12'b000001111000: finv2 = 23'b11100011010001001100100;
12'b000001111001: finv2 = 23'b11100011000010100001111;
12'b000001111010: finv2 = 23'b11100010110011110111110;
12'b000001111011: finv2 = 23'b11100010100101001110100;
12'b000001111100: finv2 = 23'b11100010010110100101110;
12'b000001111101: finv2 = 23'b11100010000111111101110;
12'b000001111110: finv2 = 23'b11100001111001010110011;
12'b000001111111: finv2 = 23'b11100001101010101111101;
12'b000010000000: finv2 = 23'b11100001011100001001101;
12'b000010000001: finv2 = 23'b11100001001101100100010;
12'b000010000010: finv2 = 23'b11100000111110111111100;
12'b000010000011: finv2 = 23'b11100000110000011011100;
12'b000010000100: finv2 = 23'b11100000100001111000001;
12'b000010000101: finv2 = 23'b11100000010011010101011;
12'b000010000110: finv2 = 23'b11100000000100110011011;
12'b000010000111: finv2 = 23'b11011111110110010010000;
12'b000010001000: finv2 = 23'b11011111100111110001010;
12'b000010001001: finv2 = 23'b11011111011001010001001;
12'b000010001010: finv2 = 23'b11011111001010110001101;
12'b000010001011: finv2 = 23'b11011110111100010010111;
12'b000010001100: finv2 = 23'b11011110101101110100110;
12'b000010001101: finv2 = 23'b11011110011111010111011;
12'b000010001110: finv2 = 23'b11011110010000111010100;
12'b000010001111: finv2 = 23'b11011110000010011110011;
12'b000010010000: finv2 = 23'b11011101110100000010111;
12'b000010010001: finv2 = 23'b11011101100101101000000;
12'b000010010010: finv2 = 23'b11011101010111001101111;
12'b000010010011: finv2 = 23'b11011101001000110100010;
12'b000010010100: finv2 = 23'b11011100111010011011011;
12'b000010010101: finv2 = 23'b11011100101100000011001;
12'b000010010110: finv2 = 23'b11011100011101101011101;
12'b000010010111: finv2 = 23'b11011100001111010100101;
12'b000010011000: finv2 = 23'b11011100000000111110011;
12'b000010011001: finv2 = 23'b11011011110010101000110;
12'b000010011010: finv2 = 23'b11011011100100010011110;
12'b000010011011: finv2 = 23'b11011011010101111111011;
12'b000010011100: finv2 = 23'b11011011000111101011101;
12'b000010011101: finv2 = 23'b11011010111001011000101;
12'b000010011110: finv2 = 23'b11011010101011000110010;
12'b000010011111: finv2 = 23'b11011010011100110100100;
12'b000010100000: finv2 = 23'b11011010001110100011011;
12'b000010100001: finv2 = 23'b11011010000000010010111;
12'b000010100010: finv2 = 23'b11011001110010000011000;
12'b000010100011: finv2 = 23'b11011001100011110011111;
12'b000010100100: finv2 = 23'b11011001010101100101010;
12'b000010100101: finv2 = 23'b11011001000111010111011;
12'b000010100110: finv2 = 23'b11011000111001001010001;
12'b000010100111: finv2 = 23'b11011000101010111101100;
12'b000010101000: finv2 = 23'b11011000011100110001100;
12'b000010101001: finv2 = 23'b11011000001110100110001;
12'b000010101010: finv2 = 23'b11011000000000011011011;
12'b000010101011: finv2 = 23'b11010111110010010001011;
12'b000010101100: finv2 = 23'b11010111100100000111111;
12'b000010101101: finv2 = 23'b11010111010101111111001;
12'b000010101110: finv2 = 23'b11010111000111110110111;
12'b000010101111: finv2 = 23'b11010110111001101111011;
12'b000010110000: finv2 = 23'b11010110101011101000100;
12'b000010110001: finv2 = 23'b11010110011101100010010;
12'b000010110010: finv2 = 23'b11010110001111011100101;
12'b000010110011: finv2 = 23'b11010110000001010111101;
12'b000010110100: finv2 = 23'b11010101110011010011010;
12'b000010110101: finv2 = 23'b11010101100101001111100;
12'b000010110110: finv2 = 23'b11010101010111001100011;
12'b000010110111: finv2 = 23'b11010101001001001001111;
12'b000010111000: finv2 = 23'b11010100111011001000001;
12'b000010111001: finv2 = 23'b11010100101101000110111;
12'b000010111010: finv2 = 23'b11010100011111000110010;
12'b000010111011: finv2 = 23'b11010100010001000110011;
12'b000010111100: finv2 = 23'b11010100000011000111000;
12'b000010111101: finv2 = 23'b11010011110101001000010;
12'b000010111110: finv2 = 23'b11010011100111001010010;
12'b000010111111: finv2 = 23'b11010011011001001100110;
12'b000011000000: finv2 = 23'b11010011001011001111111;
12'b000011000001: finv2 = 23'b11010010111101010011110;
12'b000011000010: finv2 = 23'b11010010101111011000001;
12'b000011000011: finv2 = 23'b11010010100001011101010;
12'b000011000100: finv2 = 23'b11010010010011100010111;
12'b000011000101: finv2 = 23'b11010010000101101001001;
12'b000011000110: finv2 = 23'b11010001110111110000000;
12'b000011000111: finv2 = 23'b11010001101001110111101;
12'b000011001000: finv2 = 23'b11010001011011111111110;
12'b000011001001: finv2 = 23'b11010001001110001000100;
12'b000011001010: finv2 = 23'b11010001000000010001111;
12'b000011001011: finv2 = 23'b11010000110010011011111;
12'b000011001100: finv2 = 23'b11010000100100100110100;
12'b000011001101: finv2 = 23'b11010000010110110001110;
12'b000011001110: finv2 = 23'b11010000001000111101101;
12'b000011001111: finv2 = 23'b11001111111011001010001;
12'b000011010000: finv2 = 23'b11001111101101010111010;
12'b000011010001: finv2 = 23'b11001111011111100100111;
12'b000011010010: finv2 = 23'b11001111010001110011010;
12'b000011010011: finv2 = 23'b11001111000100000010010;
12'b000011010100: finv2 = 23'b11001110110110010001110;
12'b000011010101: finv2 = 23'b11001110101000100001111;
12'b000011010110: finv2 = 23'b11001110011010110010101;
12'b000011010111: finv2 = 23'b11001110001101000100001;
12'b000011011000: finv2 = 23'b11001101111111010110001;
12'b000011011001: finv2 = 23'b11001101110001101000101;
12'b000011011010: finv2 = 23'b11001101100011111011111;
12'b000011011011: finv2 = 23'b11001101010110001111110;
12'b000011011100: finv2 = 23'b11001101001000100100001;
12'b000011011101: finv2 = 23'b11001100111010111001010;
12'b000011011110: finv2 = 23'b11001100101101001110111;
12'b000011011111: finv2 = 23'b11001100011111100101001;
12'b000011100000: finv2 = 23'b11001100010001111100000;
12'b000011100001: finv2 = 23'b11001100000100010011100;
12'b000011100010: finv2 = 23'b11001011110110101011100;
12'b000011100011: finv2 = 23'b11001011101001000100010;
12'b000011100100: finv2 = 23'b11001011011011011101100;
12'b000011100101: finv2 = 23'b11001011001101110111011;
12'b000011100110: finv2 = 23'b11001011000000010001111;
12'b000011100111: finv2 = 23'b11001010110010101101000;
12'b000011101000: finv2 = 23'b11001010100101001000110;
12'b000011101001: finv2 = 23'b11001010010111100101000;
12'b000011101010: finv2 = 23'b11001010001010000010000;
12'b000011101011: finv2 = 23'b11001001111100011111100;
12'b000011101100: finv2 = 23'b11001001101110111101100;
12'b000011101101: finv2 = 23'b11001001100001011100010;
12'b000011101110: finv2 = 23'b11001001010011111011100;
12'b000011101111: finv2 = 23'b11001001000110011011100;
12'b000011110000: finv2 = 23'b11001000111000111100000;
12'b000011110001: finv2 = 23'b11001000101011011101000;
12'b000011110010: finv2 = 23'b11001000011101111110110;
12'b000011110011: finv2 = 23'b11001000010000100001000;
12'b000011110100: finv2 = 23'b11001000000011000011111;
12'b000011110101: finv2 = 23'b11000111110101100111011;
12'b000011110110: finv2 = 23'b11000111101000001011100;
12'b000011110111: finv2 = 23'b11000111011010110000001;
12'b000011111000: finv2 = 23'b11000111001101010101011;
12'b000011111001: finv2 = 23'b11000110111111111011010;
12'b000011111010: finv2 = 23'b11000110110010100001110;
12'b000011111011: finv2 = 23'b11000110100101001000110;
12'b000011111100: finv2 = 23'b11000110010111110000011;
12'b000011111101: finv2 = 23'b11000110001010011000101;
12'b000011111110: finv2 = 23'b11000101111101000001011;
12'b000011111111: finv2 = 23'b11000101101111101010111;
12'b000100000000: finv2 = 23'b11000101100010010100111;
12'b000100000001: finv2 = 23'b11000101010100111111011;
12'b000100000010: finv2 = 23'b11000101000111101010100;
12'b000100000011: finv2 = 23'b11000100111010010110011;
12'b000100000100: finv2 = 23'b11000100101101000010101;
12'b000100000101: finv2 = 23'b11000100011111101111101;
12'b000100000110: finv2 = 23'b11000100010010011101001;
12'b000100000111: finv2 = 23'b11000100000101001011010;
12'b000100001000: finv2 = 23'b11000011110111111001111;
12'b000100001001: finv2 = 23'b11000011101010101001001;
12'b000100001010: finv2 = 23'b11000011011101011001000;
12'b000100001011: finv2 = 23'b11000011010000001001011;
12'b000100001100: finv2 = 23'b11000011000010111010100;
12'b000100001101: finv2 = 23'b11000010110101101100000;
12'b000100001110: finv2 = 23'b11000010101000011110010;
12'b000100001111: finv2 = 23'b11000010011011010001000;
12'b000100010000: finv2 = 23'b11000010001110000100011;
12'b000100010001: finv2 = 23'b11000010000000111000010;
12'b000100010010: finv2 = 23'b11000001110011101100110;
12'b000100010011: finv2 = 23'b11000001100110100001111;
12'b000100010100: finv2 = 23'b11000001011001010111100;
12'b000100010101: finv2 = 23'b11000001001100001101110;
12'b000100010110: finv2 = 23'b11000000111111000100100;
12'b000100010111: finv2 = 23'b11000000110001111011111;
12'b000100011000: finv2 = 23'b11000000100100110011111;
12'b000100011001: finv2 = 23'b11000000010111101100100;
12'b000100011010: finv2 = 23'b11000000001010100101100;
12'b000100011011: finv2 = 23'b10111111111101011111010;
12'b000100011100: finv2 = 23'b10111111110000011001100;
12'b000100011101: finv2 = 23'b10111111100011010100011;
12'b000100011110: finv2 = 23'b10111111010110001111110;
12'b000100011111: finv2 = 23'b10111111001001001011110;
12'b000100100000: finv2 = 23'b10111110111100001000010;
12'b000100100001: finv2 = 23'b10111110101111000101011;
12'b000100100010: finv2 = 23'b10111110100010000011001;
12'b000100100011: finv2 = 23'b10111110010101000001011;
12'b000100100100: finv2 = 23'b10111110001000000000010;
12'b000100100101: finv2 = 23'b10111101111010111111101;
12'b000100100110: finv2 = 23'b10111101101101111111101;
12'b000100100111: finv2 = 23'b10111101100001000000001;
12'b000100101000: finv2 = 23'b10111101010100000001010;
12'b000100101001: finv2 = 23'b10111101000111000011000;
12'b000100101010: finv2 = 23'b10111100111010000101010;
12'b000100101011: finv2 = 23'b10111100101101001000000;
12'b000100101100: finv2 = 23'b10111100100000001011011;
12'b000100101101: finv2 = 23'b10111100010011001111011;
12'b000100101110: finv2 = 23'b10111100000110010011111;
12'b000100101111: finv2 = 23'b10111011111001011001000;
12'b000100110000: finv2 = 23'b10111011101100011110101;
12'b000100110001: finv2 = 23'b10111011011111100100110;
12'b000100110010: finv2 = 23'b10111011010010101011100;
12'b000100110011: finv2 = 23'b10111011000101110010111;
12'b000100110100: finv2 = 23'b10111010111000111010110;
12'b000100110101: finv2 = 23'b10111010101100000011010;
12'b000100110110: finv2 = 23'b10111010011111001100010;
12'b000100110111: finv2 = 23'b10111010010010010101110;
12'b000100111000: finv2 = 23'b10111010000101011111111;
12'b000100111001: finv2 = 23'b10111001111000101010101;
12'b000100111010: finv2 = 23'b10111001101011110101111;
12'b000100111011: finv2 = 23'b10111001011111000001101;
12'b000100111100: finv2 = 23'b10111001010010001110000;
12'b000100111101: finv2 = 23'b10111001000101011011000;
12'b000100111110: finv2 = 23'b10111000111000101000100;
12'b000100111111: finv2 = 23'b10111000101011110110100;
12'b000101000000: finv2 = 23'b10111000011111000101001;
12'b000101000001: finv2 = 23'b10111000010010010100010;
12'b000101000010: finv2 = 23'b10111000000101100011111;
12'b000101000011: finv2 = 23'b10110111111000110100001;
12'b000101000100: finv2 = 23'b10110111101100000101000;
12'b000101000101: finv2 = 23'b10110111011111010110011;
12'b000101000110: finv2 = 23'b10110111010010101000010;
12'b000101000111: finv2 = 23'b10110111000101111010110;
12'b000101001000: finv2 = 23'b10110110111001001101110;
12'b000101001001: finv2 = 23'b10110110101100100001010;
12'b000101001010: finv2 = 23'b10110110011111110101011;
12'b000101001011: finv2 = 23'b10110110010011001010001;
12'b000101001100: finv2 = 23'b10110110000110011111010;
12'b000101001101: finv2 = 23'b10110101111001110101001;
12'b000101001110: finv2 = 23'b10110101101101001011011;
12'b000101001111: finv2 = 23'b10110101100000100010010;
12'b000101010000: finv2 = 23'b10110101010011111001101;
12'b000101010001: finv2 = 23'b10110101000111010001101;
12'b000101010010: finv2 = 23'b10110100111010101010001;
12'b000101010011: finv2 = 23'b10110100101110000011001;
12'b000101010100: finv2 = 23'b10110100100001011100110;
12'b000101010101: finv2 = 23'b10110100010100110110111;
12'b000101010110: finv2 = 23'b10110100001000010001101;
12'b000101010111: finv2 = 23'b10110011111011101100111;
12'b000101011000: finv2 = 23'b10110011101111001000101;
12'b000101011001: finv2 = 23'b10110011100010100100111;
12'b000101011010: finv2 = 23'b10110011010110000001110;
12'b000101011011: finv2 = 23'b10110011001001011111001;
12'b000101011100: finv2 = 23'b10110010111100111101001;
12'b000101011101: finv2 = 23'b10110010110000011011101;
12'b000101011110: finv2 = 23'b10110010100011111010101;
12'b000101011111: finv2 = 23'b10110010010111011010010;
12'b000101100000: finv2 = 23'b10110010001010111010011;
12'b000101100001: finv2 = 23'b10110001111110011011000;
12'b000101100010: finv2 = 23'b10110001110001111100001;
12'b000101100011: finv2 = 23'b10110001100101011101111;
12'b000101100100: finv2 = 23'b10110001011001000000001;
12'b000101100101: finv2 = 23'b10110001001100100010111;
12'b000101100110: finv2 = 23'b10110001000000000110010;
12'b000101100111: finv2 = 23'b10110000110011101010001;
12'b000101101000: finv2 = 23'b10110000100111001110100;
12'b000101101001: finv2 = 23'b10110000011010110011100;
12'b000101101010: finv2 = 23'b10110000001110011001000;
12'b000101101011: finv2 = 23'b10110000000001111111000;
12'b000101101100: finv2 = 23'b10101111110101100101100;
12'b000101101101: finv2 = 23'b10101111101001001100101;
12'b000101101110: finv2 = 23'b10101111011100110100010;
12'b000101101111: finv2 = 23'b10101111010000011100011;
12'b000101110000: finv2 = 23'b10101111000100000101000;
12'b000101110001: finv2 = 23'b10101110110111101110010;
12'b000101110010: finv2 = 23'b10101110101011011000000;
12'b000101110011: finv2 = 23'b10101110011111000010010;
12'b000101110100: finv2 = 23'b10101110010010101101001;
12'b000101110101: finv2 = 23'b10101110000110011000011;
12'b000101110110: finv2 = 23'b10101101111010000100010;
12'b000101110111: finv2 = 23'b10101101101101110000101;
12'b000101111000: finv2 = 23'b10101101100001011101101;
12'b000101111001: finv2 = 23'b10101101010101001011000;
12'b000101111010: finv2 = 23'b10101101001000111001000;
12'b000101111011: finv2 = 23'b10101100111100100111100;
12'b000101111100: finv2 = 23'b10101100110000010110100;
12'b000101111101: finv2 = 23'b10101100100100000110001;
12'b000101111110: finv2 = 23'b10101100010111110110001;
12'b000101111111: finv2 = 23'b10101100001011100110110;
12'b000110000000: finv2 = 23'b10101011111111010111111;
12'b000110000001: finv2 = 23'b10101011110011001001100;
12'b000110000010: finv2 = 23'b10101011100110111011110;
12'b000110000011: finv2 = 23'b10101011011010101110011;
12'b000110000100: finv2 = 23'b10101011001110100001101;
12'b000110000101: finv2 = 23'b10101011000010010101011;
12'b000110000110: finv2 = 23'b10101010110110001001101;
12'b000110000111: finv2 = 23'b10101010101001111110011;
12'b000110001000: finv2 = 23'b10101010011101110011110;
12'b000110001001: finv2 = 23'b10101010010001101001100;
12'b000110001010: finv2 = 23'b10101010000101011111111;
12'b000110001011: finv2 = 23'b10101001111001010110110;
12'b000110001100: finv2 = 23'b10101001101101001110001;
12'b000110001101: finv2 = 23'b10101001100001000110000;
12'b000110001110: finv2 = 23'b10101001010100111110100;
12'b000110001111: finv2 = 23'b10101001001000110111011;
12'b000110010000: finv2 = 23'b10101000111100110000111;
12'b000110010001: finv2 = 23'b10101000110000101010111;
12'b000110010010: finv2 = 23'b10101000100100100101011;
12'b000110010011: finv2 = 23'b10101000011000100000011;
12'b000110010100: finv2 = 23'b10101000001100011011111;
12'b000110010101: finv2 = 23'b10101000000000010111111;
12'b000110010110: finv2 = 23'b10100111110100010100100;
12'b000110010111: finv2 = 23'b10100111101000010001100;
12'b000110011000: finv2 = 23'b10100111011100001111001;
12'b000110011001: finv2 = 23'b10100111010000001101001;
12'b000110011010: finv2 = 23'b10100111000100001011110;
12'b000110011011: finv2 = 23'b10100110111000001010111;
12'b000110011100: finv2 = 23'b10100110101100001010100;
12'b000110011101: finv2 = 23'b10100110100000001010101;
12'b000110011110: finv2 = 23'b10100110010100001011010;
12'b000110011111: finv2 = 23'b10100110001000001100100;
12'b000110100000: finv2 = 23'b10100101111100001110001;
12'b000110100001: finv2 = 23'b10100101110000010000010;
12'b000110100010: finv2 = 23'b10100101100100010011000;
12'b000110100011: finv2 = 23'b10100101011000010110001;
12'b000110100100: finv2 = 23'b10100101001100011001111;
12'b000110100101: finv2 = 23'b10100101000000011110001;
12'b000110100110: finv2 = 23'b10100100110100100010111;
12'b000110100111: finv2 = 23'b10100100101000101000000;
12'b000110101000: finv2 = 23'b10100100011100101101110;
12'b000110101001: finv2 = 23'b10100100010000110100000;
12'b000110101010: finv2 = 23'b10100100000100111010110;
12'b000110101011: finv2 = 23'b10100011111001000010000;
12'b000110101100: finv2 = 23'b10100011101101001001110;
12'b000110101101: finv2 = 23'b10100011100001010010000;
12'b000110101110: finv2 = 23'b10100011010101011010110;
12'b000110101111: finv2 = 23'b10100011001001100100000;
12'b000110110000: finv2 = 23'b10100010111101101101110;
12'b000110110001: finv2 = 23'b10100010110001111000000;
12'b000110110010: finv2 = 23'b10100010100110000010111;
12'b000110110011: finv2 = 23'b10100010011010001110001;
12'b000110110100: finv2 = 23'b10100010001110011001111;
12'b000110110101: finv2 = 23'b10100010000010100110001;
12'b000110110110: finv2 = 23'b10100001110110110010111;
12'b000110110111: finv2 = 23'b10100001101011000000001;
12'b000110111000: finv2 = 23'b10100001011111001101111;
12'b000110111001: finv2 = 23'b10100001010011011100010;
12'b000110111010: finv2 = 23'b10100001000111101011000;
12'b000110111011: finv2 = 23'b10100000111011111010010;
12'b000110111100: finv2 = 23'b10100000110000001010000;
12'b000110111101: finv2 = 23'b10100000100100011010010;
12'b000110111110: finv2 = 23'b10100000011000101011000;
12'b000110111111: finv2 = 23'b10100000001100111100010;
12'b000111000000: finv2 = 23'b10100000000001001110000;
12'b000111000001: finv2 = 23'b10011111110101100000010;
12'b000111000010: finv2 = 23'b10011111101001110011000;
12'b000111000011: finv2 = 23'b10011111011110000110010;
12'b000111000100: finv2 = 23'b10011111010010011001111;
12'b000111000101: finv2 = 23'b10011111000110101110001;
12'b000111000110: finv2 = 23'b10011110111011000010111;
12'b000111000111: finv2 = 23'b10011110101111011000001;
12'b000111001000: finv2 = 23'b10011110100011101101110;
12'b000111001001: finv2 = 23'b10011110011000000100000;
12'b000111001010: finv2 = 23'b10011110001100011010101;
12'b000111001011: finv2 = 23'b10011110000000110001110;
12'b000111001100: finv2 = 23'b10011101110101001001100;
12'b000111001101: finv2 = 23'b10011101101001100001101;
12'b000111001110: finv2 = 23'b10011101011101111010010;
12'b000111001111: finv2 = 23'b10011101010010010011011;
12'b000111010000: finv2 = 23'b10011101000110101101000;
12'b000111010001: finv2 = 23'b10011100111011000111001;
12'b000111010010: finv2 = 23'b10011100101111100001101;
12'b000111010011: finv2 = 23'b10011100100011111100110;
12'b000111010100: finv2 = 23'b10011100011000011000011;
12'b000111010101: finv2 = 23'b10011100001100110100011;
12'b000111010110: finv2 = 23'b10011100000001010000111;
12'b000111010111: finv2 = 23'b10011011110101101110000;
12'b000111011000: finv2 = 23'b10011011101010001011100;
12'b000111011001: finv2 = 23'b10011011011110101001100;
12'b000111011010: finv2 = 23'b10011011010011001000000;
12'b000111011011: finv2 = 23'b10011011000111100110111;
12'b000111011100: finv2 = 23'b10011010111100000110011;
12'b000111011101: finv2 = 23'b10011010110000100110010;
12'b000111011110: finv2 = 23'b10011010100101000110110;
12'b000111011111: finv2 = 23'b10011010011001100111101;
12'b000111100000: finv2 = 23'b10011010001110001001000;
12'b000111100001: finv2 = 23'b10011010000010101010111;
12'b000111100010: finv2 = 23'b10011001110111001101001;
12'b000111100011: finv2 = 23'b10011001101011110000000;
12'b000111100100: finv2 = 23'b10011001100000010011010;
12'b000111100101: finv2 = 23'b10011001010100110111001;
12'b000111100110: finv2 = 23'b10011001001001011011011;
12'b000111100111: finv2 = 23'b10011000111110000000001;
12'b000111101000: finv2 = 23'b10011000110010100101010;
12'b000111101001: finv2 = 23'b10011000100111001011000;
12'b000111101010: finv2 = 23'b10011000011011110001001;
12'b000111101011: finv2 = 23'b10011000010000010111110;
12'b000111101100: finv2 = 23'b10011000000100111110111;
12'b000111101101: finv2 = 23'b10010111111001100110100;
12'b000111101110: finv2 = 23'b10010111101110001110101;
12'b000111101111: finv2 = 23'b10010111100010110111001;
12'b000111110000: finv2 = 23'b10010111010111100000010;
12'b000111110001: finv2 = 23'b10010111001100001001110;
12'b000111110010: finv2 = 23'b10010111000000110011110;
12'b000111110011: finv2 = 23'b10010110110101011110001;
12'b000111110100: finv2 = 23'b10010110101010001001001;
12'b000111110101: finv2 = 23'b10010110011110110100100;
12'b000111110110: finv2 = 23'b10010110010011100000011;
12'b000111110111: finv2 = 23'b10010110001000001100110;
12'b000111111000: finv2 = 23'b10010101111100111001100;
12'b000111111001: finv2 = 23'b10010101110001100110110;
12'b000111111010: finv2 = 23'b10010101100110010100100;
12'b000111111011: finv2 = 23'b10010101011011000010110;
12'b000111111100: finv2 = 23'b10010101001111110001100;
12'b000111111101: finv2 = 23'b10010101000100100000101;
12'b000111111110: finv2 = 23'b10010100111001010000010;
12'b000111111111: finv2 = 23'b10010100101110000000011;
12'b001000000000: finv2 = 23'b10010100100010110001000;
12'b001000000001: finv2 = 23'b10010100010111100010000;
12'b001000000010: finv2 = 23'b10010100001100010011100;
12'b001000000011: finv2 = 23'b10010100000001000101100;
12'b001000000100: finv2 = 23'b10010011110101111000000;
12'b001000000101: finv2 = 23'b10010011101010101010111;
12'b001000000110: finv2 = 23'b10010011011111011110010;
12'b001000000111: finv2 = 23'b10010011010100010010001;
12'b001000001000: finv2 = 23'b10010011001001000110011;
12'b001000001001: finv2 = 23'b10010010111101111011010;
12'b001000001010: finv2 = 23'b10010010110010110000100;
12'b001000001011: finv2 = 23'b10010010100111100110001;
12'b001000001100: finv2 = 23'b10010010011100011100011;
12'b001000001101: finv2 = 23'b10010010010001010011000;
12'b001000001110: finv2 = 23'b10010010000110001010000;
12'b001000001111: finv2 = 23'b10010001111011000001101;
12'b001000010000: finv2 = 23'b10010001101111111001101;
12'b001000010001: finv2 = 23'b10010001100100110010001;
12'b001000010010: finv2 = 23'b10010001011001101011001;
12'b001000010011: finv2 = 23'b10010001001110100100100;
12'b001000010100: finv2 = 23'b10010001000011011110011;
12'b001000010101: finv2 = 23'b10010000111000011000101;
12'b001000010110: finv2 = 23'b10010000101101010011100;
12'b001000010111: finv2 = 23'b10010000100010001110110;
12'b001000011000: finv2 = 23'b10010000010111001010011;
12'b001000011001: finv2 = 23'b10010000001100000110100;
12'b001000011010: finv2 = 23'b10010000000001000011001;
12'b001000011011: finv2 = 23'b10001111110110000000010;
12'b001000011100: finv2 = 23'b10001111101010111101110;
12'b001000011101: finv2 = 23'b10001111011111111011110;
12'b001000011110: finv2 = 23'b10001111010100111010010;
12'b001000011111: finv2 = 23'b10001111001001111001001;
12'b001000100000: finv2 = 23'b10001110111110111000100;
12'b001000100001: finv2 = 23'b10001110110011111000011;
12'b001000100010: finv2 = 23'b10001110101000111000101;
12'b001000100011: finv2 = 23'b10001110011101111001011;
12'b001000100100: finv2 = 23'b10001110010010111010100;
12'b001000100101: finv2 = 23'b10001110000111111100001;
12'b001000100110: finv2 = 23'b10001101111100111110010;
12'b001000100111: finv2 = 23'b10001101110010000000110;
12'b001000101000: finv2 = 23'b10001101100111000011110;
12'b001000101001: finv2 = 23'b10001101011100000111010;
12'b001000101010: finv2 = 23'b10001101010001001011001;
12'b001000101011: finv2 = 23'b10001101000110001111100;
12'b001000101100: finv2 = 23'b10001100111011010100010;
12'b001000101101: finv2 = 23'b10001100110000011001100;
12'b001000101110: finv2 = 23'b10001100100101011111010;
12'b001000101111: finv2 = 23'b10001100011010100101011;
12'b001000110000: finv2 = 23'b10001100001111101100000;
12'b001000110001: finv2 = 23'b10001100000100110011000;
12'b001000110010: finv2 = 23'b10001011111001111010100;
12'b001000110011: finv2 = 23'b10001011101111000010100;
12'b001000110100: finv2 = 23'b10001011100100001010111;
12'b001000110101: finv2 = 23'b10001011011001010011110;
12'b001000110110: finv2 = 23'b10001011001110011101000;
12'b001000110111: finv2 = 23'b10001011000011100110110;
12'b001000111000: finv2 = 23'b10001010111000110000111;
12'b001000111001: finv2 = 23'b10001010101101111011100;
12'b001000111010: finv2 = 23'b10001010100011000110101;
12'b001000111011: finv2 = 23'b10001010011000010010001;
12'b001000111100: finv2 = 23'b10001010001101011110001;
12'b001000111101: finv2 = 23'b10001010000010101010100;
12'b001000111110: finv2 = 23'b10001001110111110111011;
12'b001000111111: finv2 = 23'b10001001101101000100101;
12'b001001000000: finv2 = 23'b10001001100010010010011;
12'b001001000001: finv2 = 23'b10001001010111100000101;
12'b001001000010: finv2 = 23'b10001001001100101111010;
12'b001001000011: finv2 = 23'b10001001000001111110010;
12'b001001000100: finv2 = 23'b10001000110111001101111;
12'b001001000101: finv2 = 23'b10001000101100011101110;
12'b001001000110: finv2 = 23'b10001000100001101110001;
12'b001001000111: finv2 = 23'b10001000010110111111000;
12'b001001001000: finv2 = 23'b10001000001100010000010;
12'b001001001001: finv2 = 23'b10001000000001100010000;
12'b001001001010: finv2 = 23'b10000111110110110100001;
12'b001001001011: finv2 = 23'b10000111101100000110110;
12'b001001001100: finv2 = 23'b10000111100001011001110;
12'b001001001101: finv2 = 23'b10000111010110101101010;
12'b001001001110: finv2 = 23'b10000111001100000001001;
12'b001001001111: finv2 = 23'b10000111000001010101100;
12'b001001010000: finv2 = 23'b10000110110110101010011;
12'b001001010001: finv2 = 23'b10000110101011111111100;
12'b001001010010: finv2 = 23'b10000110100001010101010;
12'b001001010011: finv2 = 23'b10000110010110101011010;
12'b001001010100: finv2 = 23'b10000110001100000001111;
12'b001001010101: finv2 = 23'b10000110000001011000110;
12'b001001010110: finv2 = 23'b10000101110110110000010;
12'b001001010111: finv2 = 23'b10000101101100001000000;
12'b001001011000: finv2 = 23'b10000101100001100000011;
12'b001001011001: finv2 = 23'b10000101010110111001000;
12'b001001011010: finv2 = 23'b10000101001100010010001;
12'b001001011011: finv2 = 23'b10000101000001101011110;
12'b001001011100: finv2 = 23'b10000100110111000101110;
12'b001001011101: finv2 = 23'b10000100101100100000010;
12'b001001011110: finv2 = 23'b10000100100001111011000;
12'b001001011111: finv2 = 23'b10000100010111010110011;
12'b001001100000: finv2 = 23'b10000100001100110010001;
12'b001001100001: finv2 = 23'b10000100000010001110010;
12'b001001100010: finv2 = 23'b10000011110111101010111;
12'b001001100011: finv2 = 23'b10000011101101000111111;
12'b001001100100: finv2 = 23'b10000011100010100101011;
12'b001001100101: finv2 = 23'b10000011011000000011010;
12'b001001100110: finv2 = 23'b10000011001101100001100;
12'b001001100111: finv2 = 23'b10000011000011000000010;
12'b001001101000: finv2 = 23'b10000010111000011111100;
12'b001001101001: finv2 = 23'b10000010101101111111001;
12'b001001101010: finv2 = 23'b10000010100011011111001;
12'b001001101011: finv2 = 23'b10000010011000111111101;
12'b001001101100: finv2 = 23'b10000010001110100000100;
12'b001001101101: finv2 = 23'b10000010000100000001110;
12'b001001101110: finv2 = 23'b10000001111001100011100;
12'b001001101111: finv2 = 23'b10000001101111000101101;
12'b001001110000: finv2 = 23'b10000001100100101000010;
12'b001001110001: finv2 = 23'b10000001011010001011010;
12'b001001110010: finv2 = 23'b10000001001111101110110;
12'b001001110011: finv2 = 23'b10000001000101010010101;
12'b001001110100: finv2 = 23'b10000000111010110110111;
12'b001001110101: finv2 = 23'b10000000110000011011101;
12'b001001110110: finv2 = 23'b10000000100110000000110;
12'b001001110111: finv2 = 23'b10000000011011100110010;
12'b001001111000: finv2 = 23'b10000000010001001100010;
12'b001001111001: finv2 = 23'b10000000000110110010101;
12'b001001111010: finv2 = 23'b01111111111100011001100;
12'b001001111011: finv2 = 23'b01111111110010000000110;
12'b001001111100: finv2 = 23'b01111111100111101000011;
12'b001001111101: finv2 = 23'b01111111011101010000100;
12'b001001111110: finv2 = 23'b01111111010010111001000;
12'b001001111111: finv2 = 23'b01111111001000100010000;
12'b001010000000: finv2 = 23'b01111110111110001011011;
12'b001010000001: finv2 = 23'b01111110110011110101001;
12'b001010000010: finv2 = 23'b01111110101001011111010;
12'b001010000011: finv2 = 23'b01111110011111001001111;
12'b001010000100: finv2 = 23'b01111110010100110100111;
12'b001010000101: finv2 = 23'b01111110001010100000011;
12'b001010000110: finv2 = 23'b01111110000000001100010;
12'b001010000111: finv2 = 23'b01111101110101111000100;
12'b001010001000: finv2 = 23'b01111101101011100101010;
12'b001010001001: finv2 = 23'b01111101100001010010011;
12'b001010001010: finv2 = 23'b01111101010110111111111;
12'b001010001011: finv2 = 23'b01111101001100101101111;
12'b001010001100: finv2 = 23'b01111101000010011100001;
12'b001010001101: finv2 = 23'b01111100111000001011000;
12'b001010001110: finv2 = 23'b01111100101101111010001;
12'b001010001111: finv2 = 23'b01111100100011101001110;
12'b001010010000: finv2 = 23'b01111100011001011001110;
12'b001010010001: finv2 = 23'b01111100001111001010010;
12'b001010010010: finv2 = 23'b01111100000100111011001;
12'b001010010011: finv2 = 23'b01111011111010101100011;
12'b001010010100: finv2 = 23'b01111011110000011110000;
12'b001010010101: finv2 = 23'b01111011100110010000001;
12'b001010010110: finv2 = 23'b01111011011100000010101;
12'b001010010111: finv2 = 23'b01111011010001110101100;
12'b001010011000: finv2 = 23'b01111011000111101000111;
12'b001010011001: finv2 = 23'b01111010111101011100101;
12'b001010011010: finv2 = 23'b01111010110011010000110;
12'b001010011011: finv2 = 23'b01111010101001000101010;
12'b001010011100: finv2 = 23'b01111010011110111010010;
12'b001010011101: finv2 = 23'b01111010010100101111101;
12'b001010011110: finv2 = 23'b01111010001010100101100;
12'b001010011111: finv2 = 23'b01111010000000011011101;
12'b001010100000: finv2 = 23'b01111001110110010010010;
12'b001010100001: finv2 = 23'b01111001101100001001010;
12'b001010100010: finv2 = 23'b01111001100010000000101;
12'b001010100011: finv2 = 23'b01111001010111111000100;
12'b001010100100: finv2 = 23'b01111001001101110000110;
12'b001010100101: finv2 = 23'b01111001000011101001011;
12'b001010100110: finv2 = 23'b01111000111001100010100;
12'b001010100111: finv2 = 23'b01111000101111011011111;
12'b001010101000: finv2 = 23'b01111000100101010101110;
12'b001010101001: finv2 = 23'b01111000011011010000000;
12'b001010101010: finv2 = 23'b01111000010001001010110;
12'b001010101011: finv2 = 23'b01111000000111000101110;
12'b001010101100: finv2 = 23'b01110111111101000001010;
12'b001010101101: finv2 = 23'b01110111110010111101001;
12'b001010101110: finv2 = 23'b01110111101000111001100;
12'b001010101111: finv2 = 23'b01110111011110110110001;
12'b001010110000: finv2 = 23'b01110111010100110011010;
12'b001010110001: finv2 = 23'b01110111001010110000110;
12'b001010110010: finv2 = 23'b01110111000000101110110;
12'b001010110011: finv2 = 23'b01110110110110101101000;
12'b001010110100: finv2 = 23'b01110110101100101011110;
12'b001010110101: finv2 = 23'b01110110100010101010111;
12'b001010110110: finv2 = 23'b01110110011000101010011;
12'b001010110111: finv2 = 23'b01110110001110101010010;
12'b001010111000: finv2 = 23'b01110110000100101010101;
12'b001010111001: finv2 = 23'b01110101111010101011010;
12'b001010111010: finv2 = 23'b01110101110000101100011;
12'b001010111011: finv2 = 23'b01110101100110101101111;
12'b001010111100: finv2 = 23'b01110101011100101111111;
12'b001010111101: finv2 = 23'b01110101010010110010001;
12'b001010111110: finv2 = 23'b01110101001000110100111;
12'b001010111111: finv2 = 23'b01110100111110111000000;
12'b001011000000: finv2 = 23'b01110100110100111011100;
12'b001011000001: finv2 = 23'b01110100101010111111011;
12'b001011000010: finv2 = 23'b01110100100001000011110;
12'b001011000011: finv2 = 23'b01110100010111001000011;
12'b001011000100: finv2 = 23'b01110100001101001101100;
12'b001011000101: finv2 = 23'b01110100000011010011000;
12'b001011000110: finv2 = 23'b01110011111001011000111;
12'b001011000111: finv2 = 23'b01110011101111011111001;
12'b001011001000: finv2 = 23'b01110011100101100101111;
12'b001011001001: finv2 = 23'b01110011011011101100111;
12'b001011001010: finv2 = 23'b01110011010001110100011;
12'b001011001011: finv2 = 23'b01110011000111111100010;
12'b001011001100: finv2 = 23'b01110010111110000100100;
12'b001011001101: finv2 = 23'b01110010110100001101001;
12'b001011001110: finv2 = 23'b01110010101010010110010;
12'b001011001111: finv2 = 23'b01110010100000011111101;
12'b001011010000: finv2 = 23'b01110010010110101001100;
12'b001011010001: finv2 = 23'b01110010001100110011110;
12'b001011010010: finv2 = 23'b01110010000010111110011;
12'b001011010011: finv2 = 23'b01110001111001001001011;
12'b001011010100: finv2 = 23'b01110001101111010100110;
12'b001011010101: finv2 = 23'b01110001100101100000100;
12'b001011010110: finv2 = 23'b01110001011011101100110;
12'b001011010111: finv2 = 23'b01110001010001111001010;
12'b001011011000: finv2 = 23'b01110001001000000110010;
12'b001011011001: finv2 = 23'b01110000111110010011101;
12'b001011011010: finv2 = 23'b01110000110100100001011;
12'b001011011011: finv2 = 23'b01110000101010101111100;
12'b001011011100: finv2 = 23'b01110000100000111110000;
12'b001011011101: finv2 = 23'b01110000010111001100111;
12'b001011011110: finv2 = 23'b01110000001101011100010;
12'b001011011111: finv2 = 23'b01110000000011101011111;
12'b001011100000: finv2 = 23'b01101111111001111100000;
12'b001011100001: finv2 = 23'b01101111110000001100011;
12'b001011100010: finv2 = 23'b01101111100110011101010;
12'b001011100011: finv2 = 23'b01101111011100101110100;
12'b001011100100: finv2 = 23'b01101111010011000000001;
12'b001011100101: finv2 = 23'b01101111001001010010001;
12'b001011100110: finv2 = 23'b01101110111111100100100;
12'b001011100111: finv2 = 23'b01101110110101110111010;
12'b001011101000: finv2 = 23'b01101110101100001010100;
12'b001011101001: finv2 = 23'b01101110100010011110000;
12'b001011101010: finv2 = 23'b01101110011000110010000;
12'b001011101011: finv2 = 23'b01101110001111000110010;
12'b001011101100: finv2 = 23'b01101110000101011011000;
12'b001011101101: finv2 = 23'b01101101111011110000000;
12'b001011101110: finv2 = 23'b01101101110010000101100;
12'b001011101111: finv2 = 23'b01101101101000011011011;
12'b001011110000: finv2 = 23'b01101101011110110001101;
12'b001011110001: finv2 = 23'b01101101010101001000010;
12'b001011110010: finv2 = 23'b01101101001011011111010;
12'b001011110011: finv2 = 23'b01101101000001110110101;
12'b001011110100: finv2 = 23'b01101100111000001110011;
12'b001011110101: finv2 = 23'b01101100101110100110100;
12'b001011110110: finv2 = 23'b01101100100100111111000;
12'b001011110111: finv2 = 23'b01101100011011010111111;
12'b001011111000: finv2 = 23'b01101100010001110001001;
12'b001011111001: finv2 = 23'b01101100001000001010111;
12'b001011111010: finv2 = 23'b01101011111110100100111;
12'b001011111011: finv2 = 23'b01101011110100111111010;
12'b001011111100: finv2 = 23'b01101011101011011010001;
12'b001011111101: finv2 = 23'b01101011100001110101010;
12'b001011111110: finv2 = 23'b01101011011000010000110;
12'b001011111111: finv2 = 23'b01101011001110101100110;
12'b001100000000: finv2 = 23'b01101011000101001001000;
12'b001100000001: finv2 = 23'b01101010111011100101110;
12'b001100000010: finv2 = 23'b01101010110010000010110;
12'b001100000011: finv2 = 23'b01101010101000100000010;
12'b001100000100: finv2 = 23'b01101010011110111110000;
12'b001100000101: finv2 = 23'b01101010010101011100010;
12'b001100000110: finv2 = 23'b01101010001011111010110;
12'b001100000111: finv2 = 23'b01101010000010011001110;
12'b001100001000: finv2 = 23'b01101001111000111001000;
12'b001100001001: finv2 = 23'b01101001101111011000110;
12'b001100001010: finv2 = 23'b01101001100101111000110;
12'b001100001011: finv2 = 23'b01101001011100011001010;
12'b001100001100: finv2 = 23'b01101001010010111010001;
12'b001100001101: finv2 = 23'b01101001001001011011010;
12'b001100001110: finv2 = 23'b01101000111111111100110;
12'b001100001111: finv2 = 23'b01101000110110011110110;
12'b001100010000: finv2 = 23'b01101000101101000001000;
12'b001100010001: finv2 = 23'b01101000100011100011110;
12'b001100010010: finv2 = 23'b01101000011010000110110;
12'b001100010011: finv2 = 23'b01101000010000101010010;
12'b001100010100: finv2 = 23'b01101000000111001110000;
12'b001100010101: finv2 = 23'b01100111111101110010001;
12'b001100010110: finv2 = 23'b01100111110100010110101;
12'b001100010111: finv2 = 23'b01100111101010111011101;
12'b001100011000: finv2 = 23'b01100111100001100000111;
12'b001100011001: finv2 = 23'b01100111011000000110100;
12'b001100011010: finv2 = 23'b01100111001110101100100;
12'b001100011011: finv2 = 23'b01100111000101010010111;
12'b001100011100: finv2 = 23'b01100110111011111001101;
12'b001100011101: finv2 = 23'b01100110110010100000110;
12'b001100011110: finv2 = 23'b01100110101001001000010;
12'b001100011111: finv2 = 23'b01100110011111110000001;
12'b001100100000: finv2 = 23'b01100110010110011000011;
12'b001100100001: finv2 = 23'b01100110001101000001000;
12'b001100100010: finv2 = 23'b01100110000011101001111;
12'b001100100011: finv2 = 23'b01100101111010010011010;
12'b001100100100: finv2 = 23'b01100101110000111100111;
12'b001100100101: finv2 = 23'b01100101100111100111000;
12'b001100100110: finv2 = 23'b01100101011110010001011;
12'b001100100111: finv2 = 23'b01100101010100111100010;
12'b001100101000: finv2 = 23'b01100101001011100111011;
12'b001100101001: finv2 = 23'b01100101000010010010111;
12'b001100101010: finv2 = 23'b01100100111000111110110;
12'b001100101011: finv2 = 23'b01100100101111101011000;
12'b001100101100: finv2 = 23'b01100100100110010111101;
12'b001100101101: finv2 = 23'b01100100011101000100101;
12'b001100101110: finv2 = 23'b01100100010011110001111;
12'b001100101111: finv2 = 23'b01100100001010011111101;
12'b001100110000: finv2 = 23'b01100100000001001101110;
12'b001100110001: finv2 = 23'b01100011110111111100001;
12'b001100110010: finv2 = 23'b01100011101110101010111;
12'b001100110011: finv2 = 23'b01100011100101011010001;
12'b001100110100: finv2 = 23'b01100011011100001001101;
12'b001100110101: finv2 = 23'b01100011010010111001100;
12'b001100110110: finv2 = 23'b01100011001001101001110;
12'b001100110111: finv2 = 23'b01100011000000011010010;
12'b001100111000: finv2 = 23'b01100010110111001011010;
12'b001100111001: finv2 = 23'b01100010101101111100101;
12'b001100111010: finv2 = 23'b01100010100100101110010;
12'b001100111011: finv2 = 23'b01100010011011100000011;
12'b001100111100: finv2 = 23'b01100010010010010010110;
12'b001100111101: finv2 = 23'b01100010001001000101100;
12'b001100111110: finv2 = 23'b01100001111111111000101;
12'b001100111111: finv2 = 23'b01100001110110101100001;
12'b001101000000: finv2 = 23'b01100001101101011111111;
12'b001101000001: finv2 = 23'b01100001100100010100001;
12'b001101000010: finv2 = 23'b01100001011011001000101;
12'b001101000011: finv2 = 23'b01100001010001111101100;
12'b001101000100: finv2 = 23'b01100001001000110010110;
12'b001101000101: finv2 = 23'b01100000111111101000011;
12'b001101000110: finv2 = 23'b01100000110110011110011;
12'b001101000111: finv2 = 23'b01100000101101010100110;
12'b001101001000: finv2 = 23'b01100000100100001011011;
12'b001101001001: finv2 = 23'b01100000011011000010100;
12'b001101001010: finv2 = 23'b01100000010001111001111;
12'b001101001011: finv2 = 23'b01100000001000110001101;
12'b001101001100: finv2 = 23'b01011111111111101001110;
12'b001101001101: finv2 = 23'b01011111110110100010010;
12'b001101001110: finv2 = 23'b01011111101101011011000;
12'b001101001111: finv2 = 23'b01011111100100010100010;
12'b001101010000: finv2 = 23'b01011111011011001101110;
12'b001101010001: finv2 = 23'b01011111010010000111101;
12'b001101010010: finv2 = 23'b01011111001001000001111;
12'b001101010011: finv2 = 23'b01011110111111111100011;
12'b001101010100: finv2 = 23'b01011110110110110111011;
12'b001101010101: finv2 = 23'b01011110101101110010101;
12'b001101010110: finv2 = 23'b01011110100100101110010;
12'b001101010111: finv2 = 23'b01011110011011101010010;
12'b001101011000: finv2 = 23'b01011110010010100110101;
12'b001101011001: finv2 = 23'b01011110001001100011011;
12'b001101011010: finv2 = 23'b01011110000000100000011;
12'b001101011011: finv2 = 23'b01011101110111011101110;
12'b001101011100: finv2 = 23'b01011101101110011011100;
12'b001101011101: finv2 = 23'b01011101100101011001101;
12'b001101011110: finv2 = 23'b01011101011100011000001;
12'b001101011111: finv2 = 23'b01011101010011010110111;
12'b001101100000: finv2 = 23'b01011101001010010110000;
12'b001101100001: finv2 = 23'b01011101000001010101100;
12'b001101100010: finv2 = 23'b01011100111000010101011;
12'b001101100011: finv2 = 23'b01011100101111010101100;
12'b001101100100: finv2 = 23'b01011100100110010110001;
12'b001101100101: finv2 = 23'b01011100011101010111000;
12'b001101100110: finv2 = 23'b01011100010100011000010;
12'b001101100111: finv2 = 23'b01011100001011011001110;
12'b001101101000: finv2 = 23'b01011100000010011011110;
12'b001101101001: finv2 = 23'b01011011111001011110000;
12'b001101101010: finv2 = 23'b01011011110000100000101;
12'b001101101011: finv2 = 23'b01011011100111100011101;
12'b001101101100: finv2 = 23'b01011011011110100110111;
12'b001101101101: finv2 = 23'b01011011010101101010100;
12'b001101101110: finv2 = 23'b01011011001100101110100;
12'b001101101111: finv2 = 23'b01011011000011110010111;
12'b001101110000: finv2 = 23'b01011010111010110111101;
12'b001101110001: finv2 = 23'b01011010110001111100101;
12'b001101110010: finv2 = 23'b01011010101001000010000;
12'b001101110011: finv2 = 23'b01011010100000000111110;
12'b001101110100: finv2 = 23'b01011010010111001101110;
12'b001101110101: finv2 = 23'b01011010001110010100010;
12'b001101110110: finv2 = 23'b01011010000101011011000;
12'b001101110111: finv2 = 23'b01011001111100100010001;
12'b001101111000: finv2 = 23'b01011001110011101001100;
12'b001101111001: finv2 = 23'b01011001101010110001010;
12'b001101111010: finv2 = 23'b01011001100001111001011;
12'b001101111011: finv2 = 23'b01011001011001000001111;
12'b001101111100: finv2 = 23'b01011001010000001010101;
12'b001101111101: finv2 = 23'b01011001000111010011111;
12'b001101111110: finv2 = 23'b01011000111110011101011;
12'b001101111111: finv2 = 23'b01011000110101100111001;
12'b001110000000: finv2 = 23'b01011000101100110001011;
12'b001110000001: finv2 = 23'b01011000100011111011111;
12'b001110000010: finv2 = 23'b01011000011011000110101;
12'b001110000011: finv2 = 23'b01011000010010010001111;
12'b001110000100: finv2 = 23'b01011000001001011101011;
12'b001110000101: finv2 = 23'b01011000000000101001010;
12'b001110000110: finv2 = 23'b01010111110111110101100;
12'b001110000111: finv2 = 23'b01010111101111000010000;
12'b001110001000: finv2 = 23'b01010111100110001110111;
12'b001110001001: finv2 = 23'b01010111011101011100001;
12'b001110001010: finv2 = 23'b01010111010100101001101;
12'b001110001011: finv2 = 23'b01010111001011110111100;
12'b001110001100: finv2 = 23'b01010111000011000101110;
12'b001110001101: finv2 = 23'b01010110111010010100011;
12'b001110001110: finv2 = 23'b01010110110001100011010;
12'b001110001111: finv2 = 23'b01010110101000110010100;
12'b001110010000: finv2 = 23'b01010110100000000010001;
12'b001110010001: finv2 = 23'b01010110010111010010000;
12'b001110010010: finv2 = 23'b01010110001110100010010;
12'b001110010011: finv2 = 23'b01010110000101110010110;
12'b001110010100: finv2 = 23'b01010101111101000011110;
12'b001110010101: finv2 = 23'b01010101110100010101000;
12'b001110010110: finv2 = 23'b01010101101011100110101;
12'b001110010111: finv2 = 23'b01010101100010111000100;
12'b001110011000: finv2 = 23'b01010101011010001010110;
12'b001110011001: finv2 = 23'b01010101010001011101011;
12'b001110011010: finv2 = 23'b01010101001000110000010;
12'b001110011011: finv2 = 23'b01010101000000000011100;
12'b001110011100: finv2 = 23'b01010100110111010111001;
12'b001110011101: finv2 = 23'b01010100101110101011000;
12'b001110011110: finv2 = 23'b01010100100101111111010;
12'b001110011111: finv2 = 23'b01010100011101010011111;
12'b001110100000: finv2 = 23'b01010100010100101000110;
12'b001110100001: finv2 = 23'b01010100001011111110000;
12'b001110100010: finv2 = 23'b01010100000011010011101;
12'b001110100011: finv2 = 23'b01010011111010101001100;
12'b001110100100: finv2 = 23'b01010011110001111111110;
12'b001110100101: finv2 = 23'b01010011101001010110010;
12'b001110100110: finv2 = 23'b01010011100000101101001;
12'b001110100111: finv2 = 23'b01010011011000000100011;
12'b001110101000: finv2 = 23'b01010011001111011100000;
12'b001110101001: finv2 = 23'b01010011000110110011111;
12'b001110101010: finv2 = 23'b01010010111110001100000;
12'b001110101011: finv2 = 23'b01010010110101100100101;
12'b001110101100: finv2 = 23'b01010010101100111101100;
12'b001110101101: finv2 = 23'b01010010100100010110101;
12'b001110101110: finv2 = 23'b01010010011011110000010;
12'b001110101111: finv2 = 23'b01010010010011001010001;
12'b001110110000: finv2 = 23'b01010010001010100100010;
12'b001110110001: finv2 = 23'b01010010000001111110110;
12'b001110110010: finv2 = 23'b01010001111001011001101;
12'b001110110011: finv2 = 23'b01010001110000110100110;
12'b001110110100: finv2 = 23'b01010001101000010000010;
12'b001110110101: finv2 = 23'b01010001011111101100001;
12'b001110110110: finv2 = 23'b01010001010111001000010;
12'b001110110111: finv2 = 23'b01010001001110100100101;
12'b001110111000: finv2 = 23'b01010001000110000001100;
12'b001110111001: finv2 = 23'b01010000111101011110101;
12'b001110111010: finv2 = 23'b01010000110100111100000;
12'b001110111011: finv2 = 23'b01010000101100011001110;
12'b001110111100: finv2 = 23'b01010000100011110111111;
12'b001110111101: finv2 = 23'b01010000011011010110011;
12'b001110111110: finv2 = 23'b01010000010010110101000;
12'b001110111111: finv2 = 23'b01010000001010010100001;
12'b001111000000: finv2 = 23'b01010000000001110011100;
12'b001111000001: finv2 = 23'b01001111111001010011010;
12'b001111000010: finv2 = 23'b01001111110000110011010;
12'b001111000011: finv2 = 23'b01001111101000010011101;
12'b001111000100: finv2 = 23'b01001111011111110100010;
12'b001111000101: finv2 = 23'b01001111010111010101010;
12'b001111000110: finv2 = 23'b01001111001110110110101;
12'b001111000111: finv2 = 23'b01001111000110011000010;
12'b001111001000: finv2 = 23'b01001110111101111010010;
12'b001111001001: finv2 = 23'b01001110110101011100100;
12'b001111001010: finv2 = 23'b01001110101100111111001;
12'b001111001011: finv2 = 23'b01001110100100100010000;
12'b001111001100: finv2 = 23'b01001110011100000101010;
12'b001111001101: finv2 = 23'b01001110010011101000111;
12'b001111001110: finv2 = 23'b01001110001011001100110;
12'b001111001111: finv2 = 23'b01001110000010110001000;
12'b001111010000: finv2 = 23'b01001101111010010101100;
12'b001111010001: finv2 = 23'b01001101110001111010011;
12'b001111010010: finv2 = 23'b01001101101001011111100;
12'b001111010011: finv2 = 23'b01001101100001000101000;
12'b001111010100: finv2 = 23'b01001101011000101010110;
12'b001111010101: finv2 = 23'b01001101010000010000111;
12'b001111010110: finv2 = 23'b01001101000111110111011;
12'b001111010111: finv2 = 23'b01001100111111011110001;
12'b001111011000: finv2 = 23'b01001100110111000101001;
12'b001111011001: finv2 = 23'b01001100101110101100100;
12'b001111011010: finv2 = 23'b01001100100110010100010;
12'b001111011011: finv2 = 23'b01001100011101111100010;
12'b001111011100: finv2 = 23'b01001100010101100100101;
12'b001111011101: finv2 = 23'b01001100001101001101010;
12'b001111011110: finv2 = 23'b01001100000100110110010;
12'b001111011111: finv2 = 23'b01001011111100011111100;
12'b001111100000: finv2 = 23'b01001011110100001001001;
12'b001111100001: finv2 = 23'b01001011101011110011000;
12'b001111100010: finv2 = 23'b01001011100011011101010;
12'b001111100011: finv2 = 23'b01001011011011000111110;
12'b001111100100: finv2 = 23'b01001011010010110010101;
12'b001111100101: finv2 = 23'b01001011001010011101111;
12'b001111100110: finv2 = 23'b01001011000010001001010;
12'b001111100111: finv2 = 23'b01001010111001110101001;
12'b001111101000: finv2 = 23'b01001010110001100001010;
12'b001111101001: finv2 = 23'b01001010101001001101101;
12'b001111101010: finv2 = 23'b01001010100000111010011;
12'b001111101011: finv2 = 23'b01001010011000100111100;
12'b001111101100: finv2 = 23'b01001010010000010100110;
12'b001111101101: finv2 = 23'b01001010001000000010100;
12'b001111101110: finv2 = 23'b01001001111111110000100;
12'b001111101111: finv2 = 23'b01001001110111011110110;
12'b001111110000: finv2 = 23'b01001001101111001101011;
12'b001111110001: finv2 = 23'b01001001100110111100010;
12'b001111110010: finv2 = 23'b01001001011110101011100;
12'b001111110011: finv2 = 23'b01001001010110011011001;
12'b001111110100: finv2 = 23'b01001001001110001010111;
12'b001111110101: finv2 = 23'b01001001000101111011001;
12'b001111110110: finv2 = 23'b01001000111101101011100;
12'b001111110111: finv2 = 23'b01001000110101011100011;
12'b001111111000: finv2 = 23'b01001000101101001101011;
12'b001111111001: finv2 = 23'b01001000100100111110111;
12'b001111111010: finv2 = 23'b01001000011100110000100;
12'b001111111011: finv2 = 23'b01001000010100100010101;
12'b001111111100: finv2 = 23'b01001000001100010100111;
12'b001111111101: finv2 = 23'b01001000000100000111100;
12'b001111111110: finv2 = 23'b01000111111011111010100;
12'b001111111111: finv2 = 23'b01000111110011101101110;
12'b010000000000: finv2 = 23'b01000111101011100001010;
12'b010000000001: finv2 = 23'b01000111100011010101001;
12'b010000000010: finv2 = 23'b01000111011011001001011;
12'b010000000011: finv2 = 23'b01000111010010111101110;
12'b010000000100: finv2 = 23'b01000111001010110010101;
12'b010000000101: finv2 = 23'b01000111000010100111101;
12'b010000000110: finv2 = 23'b01000110111010011101001;
12'b010000000111: finv2 = 23'b01000110110010010010110;
12'b010000001000: finv2 = 23'b01000110101010001000110;
12'b010000001001: finv2 = 23'b01000110100001111111001;
12'b010000001010: finv2 = 23'b01000110011001110101110;
12'b010000001011: finv2 = 23'b01000110010001101100101;
12'b010000001100: finv2 = 23'b01000110001001100011111;
12'b010000001101: finv2 = 23'b01000110000001011011011;
12'b010000001110: finv2 = 23'b01000101111001010011010;
12'b010000001111: finv2 = 23'b01000101110001001011011;
12'b010000010000: finv2 = 23'b01000101101001000011111;
12'b010000010001: finv2 = 23'b01000101100000111100101;
12'b010000010010: finv2 = 23'b01000101011000110101101;
12'b010000010011: finv2 = 23'b01000101010000101111000;
12'b010000010100: finv2 = 23'b01000101001000101000101;
12'b010000010101: finv2 = 23'b01000101000000100010101;
12'b010000010110: finv2 = 23'b01000100111000011100111;
12'b010000010111: finv2 = 23'b01000100110000010111011;
12'b010000011000: finv2 = 23'b01000100101000010010010;
12'b010000011001: finv2 = 23'b01000100100000001101100;
12'b010000011010: finv2 = 23'b01000100011000001000111;
12'b010000011011: finv2 = 23'b01000100010000000100110;
12'b010000011100: finv2 = 23'b01000100001000000000110;
12'b010000011101: finv2 = 23'b01000011111111111101001;
12'b010000011110: finv2 = 23'b01000011110111111001110;
12'b010000011111: finv2 = 23'b01000011101111110110110;
12'b010000100000: finv2 = 23'b01000011100111110100000;
12'b010000100001: finv2 = 23'b01000011011111110001101;
12'b010000100010: finv2 = 23'b01000011010111101111100;
12'b010000100011: finv2 = 23'b01000011001111101101101;
12'b010000100100: finv2 = 23'b01000011000111101100001;
12'b010000100101: finv2 = 23'b01000010111111101010111;
12'b010000100110: finv2 = 23'b01000010110111101010000;
12'b010000100111: finv2 = 23'b01000010101111101001011;
12'b010000101000: finv2 = 23'b01000010100111101001000;
12'b010000101001: finv2 = 23'b01000010011111101001000;
12'b010000101010: finv2 = 23'b01000010010111101001010;
12'b010000101011: finv2 = 23'b01000010001111101001110;
12'b010000101100: finv2 = 23'b01000010000111101010101;
12'b010000101101: finv2 = 23'b01000001111111101011110;
12'b010000101110: finv2 = 23'b01000001110111101101010;
12'b010000101111: finv2 = 23'b01000001101111101111000;
12'b010000110000: finv2 = 23'b01000001100111110001000;
12'b010000110001: finv2 = 23'b01000001011111110011010;
12'b010000110010: finv2 = 23'b01000001010111110110000;
12'b010000110011: finv2 = 23'b01000001001111111000111;
12'b010000110100: finv2 = 23'b01000001000111111100001;
12'b010000110101: finv2 = 23'b01000000111111111111101;
12'b010000110110: finv2 = 23'b01000000111000000011011;
12'b010000110111: finv2 = 23'b01000000110000000111100;
12'b010000111000: finv2 = 23'b01000000101000001011111;
12'b010000111001: finv2 = 23'b01000000100000010000101;
12'b010000111010: finv2 = 23'b01000000011000010101101;
12'b010000111011: finv2 = 23'b01000000010000011010111;
12'b010000111100: finv2 = 23'b01000000001000100000100;
12'b010000111101: finv2 = 23'b01000000000000100110010;
12'b010000111110: finv2 = 23'b00111111111000101100100;
12'b010000111111: finv2 = 23'b00111111110000110010111;
12'b010001000000: finv2 = 23'b00111111101000111001101;
12'b010001000001: finv2 = 23'b00111111100001000000110;
12'b010001000010: finv2 = 23'b00111111011001001000000;
12'b010001000011: finv2 = 23'b00111111010001001111101;
12'b010001000100: finv2 = 23'b00111111001001010111101;
12'b010001000101: finv2 = 23'b00111111000001011111110;
12'b010001000110: finv2 = 23'b00111110111001101000010;
12'b010001000111: finv2 = 23'b00111110110001110001000;
12'b010001001000: finv2 = 23'b00111110101001111010001;
12'b010001001001: finv2 = 23'b00111110100010000011100;
12'b010001001010: finv2 = 23'b00111110011010001101001;
12'b010001001011: finv2 = 23'b00111110010010010111001;
12'b010001001100: finv2 = 23'b00111110001010100001011;
12'b010001001101: finv2 = 23'b00111110000010101011111;
12'b010001001110: finv2 = 23'b00111101111010110110110;
12'b010001001111: finv2 = 23'b00111101110011000001110;
12'b010001010000: finv2 = 23'b00111101101011001101010;
12'b010001010001: finv2 = 23'b00111101100011011000111;
12'b010001010010: finv2 = 23'b00111101011011100100111;
12'b010001010011: finv2 = 23'b00111101010011110001001;
12'b010001010100: finv2 = 23'b00111101001011111101101;
12'b010001010101: finv2 = 23'b00111101000100001010100;
12'b010001010110: finv2 = 23'b00111100111100010111101;
12'b010001010111: finv2 = 23'b00111100110100100101000;
12'b010001011000: finv2 = 23'b00111100101100110010110;
12'b010001011001: finv2 = 23'b00111100100101000000110;
12'b010001011010: finv2 = 23'b00111100011101001111000;
12'b010001011011: finv2 = 23'b00111100010101011101100;
12'b010001011100: finv2 = 23'b00111100001101101100011;
12'b010001011101: finv2 = 23'b00111100000101111011100;
12'b010001011110: finv2 = 23'b00111011111110001011000;
12'b010001011111: finv2 = 23'b00111011110110011010101;
12'b010001100000: finv2 = 23'b00111011101110101010101;
12'b010001100001: finv2 = 23'b00111011100110111010111;
12'b010001100010: finv2 = 23'b00111011011111001011100;
12'b010001100011: finv2 = 23'b00111011010111011100010;
12'b010001100100: finv2 = 23'b00111011001111101101011;
12'b010001100101: finv2 = 23'b00111011000111111110111;
12'b010001100110: finv2 = 23'b00111011000000010000100;
12'b010001100111: finv2 = 23'b00111010111000100010100;
12'b010001101000: finv2 = 23'b00111010110000110100110;
12'b010001101001: finv2 = 23'b00111010101001000111011;
12'b010001101010: finv2 = 23'b00111010100001011010001;
12'b010001101011: finv2 = 23'b00111010011001101101010;
12'b010001101100: finv2 = 23'b00111010010010000000101;
12'b010001101101: finv2 = 23'b00111010001010010100011;
12'b010001101110: finv2 = 23'b00111010000010101000011;
12'b010001101111: finv2 = 23'b00111001111010111100100;
12'b010001110000: finv2 = 23'b00111001110011010001001;
12'b010001110001: finv2 = 23'b00111001101011100101111;
12'b010001110010: finv2 = 23'b00111001100011111011000;
12'b010001110011: finv2 = 23'b00111001011100010000011;
12'b010001110100: finv2 = 23'b00111001010100100110000;
12'b010001110101: finv2 = 23'b00111001001100111011111;
12'b010001110110: finv2 = 23'b00111001000101010010001;
12'b010001110111: finv2 = 23'b00111000111101101000101;
12'b010001111000: finv2 = 23'b00111000110101111111011;
12'b010001111001: finv2 = 23'b00111000101110010110100;
12'b010001111010: finv2 = 23'b00111000100110101101110;
12'b010001111011: finv2 = 23'b00111000011111000101011;
12'b010001111100: finv2 = 23'b00111000010111011101010;
12'b010001111101: finv2 = 23'b00111000001111110101100;
12'b010001111110: finv2 = 23'b00111000001000001101111;
12'b010001111111: finv2 = 23'b00111000000000100110101;
12'b010010000000: finv2 = 23'b00110111111000111111101;
12'b010010000001: finv2 = 23'b00110111110001011001000;
12'b010010000010: finv2 = 23'b00110111101001110010100;
12'b010010000011: finv2 = 23'b00110111100010001100011;
12'b010010000100: finv2 = 23'b00110111011010100110100;
12'b010010000101: finv2 = 23'b00110111010011000000111;
12'b010010000110: finv2 = 23'b00110111001011011011100;
12'b010010000111: finv2 = 23'b00110111000011110110100;
12'b010010001000: finv2 = 23'b00110110111100010001110;
12'b010010001001: finv2 = 23'b00110110110100101101010;
12'b010010001010: finv2 = 23'b00110110101101001001000;
12'b010010001011: finv2 = 23'b00110110100101100101000;
12'b010010001100: finv2 = 23'b00110110011110000001011;
12'b010010001101: finv2 = 23'b00110110010110011110000;
12'b010010001110: finv2 = 23'b00110110001110111010111;
12'b010010001111: finv2 = 23'b00110110000111011000000;
12'b010010010000: finv2 = 23'b00110101111111110101100;
12'b010010010001: finv2 = 23'b00110101111000010011010;
12'b010010010010: finv2 = 23'b00110101110000110001001;
12'b010010010011: finv2 = 23'b00110101101001001111011;
12'b010010010100: finv2 = 23'b00110101100001101110000;
12'b010010010101: finv2 = 23'b00110101011010001100110;
12'b010010010110: finv2 = 23'b00110101010010101011111;
12'b010010010111: finv2 = 23'b00110101001011001011010;
12'b010010011000: finv2 = 23'b00110101000011101010111;
12'b010010011001: finv2 = 23'b00110100111100001010110;
12'b010010011010: finv2 = 23'b00110100110100101010111;
12'b010010011011: finv2 = 23'b00110100101101001011011;
12'b010010011100: finv2 = 23'b00110100100101101100001;
12'b010010011101: finv2 = 23'b00110100011110001101001;
12'b010010011110: finv2 = 23'b00110100010110101110011;
12'b010010011111: finv2 = 23'b00110100001111001111111;
12'b010010100000: finv2 = 23'b00110100000111110001110;
12'b010010100001: finv2 = 23'b00110100000000010011110;
12'b010010100010: finv2 = 23'b00110011111000110110001;
12'b010010100011: finv2 = 23'b00110011110001011000110;
12'b010010100100: finv2 = 23'b00110011101001111011101;
12'b010010100101: finv2 = 23'b00110011100010011110110;
12'b010010100110: finv2 = 23'b00110011011011000010010;
12'b010010100111: finv2 = 23'b00110011010011100110000;
12'b010010101000: finv2 = 23'b00110011001100001001111;
12'b010010101001: finv2 = 23'b00110011000100101110001;
12'b010010101010: finv2 = 23'b00110010111101010010101;
12'b010010101011: finv2 = 23'b00110010110101110111100;
12'b010010101100: finv2 = 23'b00110010101110011100100;
12'b010010101101: finv2 = 23'b00110010100111000001111;
12'b010010101110: finv2 = 23'b00110010011111100111100;
12'b010010101111: finv2 = 23'b00110010011000001101010;
12'b010010110000: finv2 = 23'b00110010010000110011011;
12'b010010110001: finv2 = 23'b00110010001001011001111;
12'b010010110010: finv2 = 23'b00110010000010000000100;
12'b010010110011: finv2 = 23'b00110001111010100111011;
12'b010010110100: finv2 = 23'b00110001110011001110101;
12'b010010110101: finv2 = 23'b00110001101011110110001;
12'b010010110110: finv2 = 23'b00110001100100011101111;
12'b010010110111: finv2 = 23'b00110001011101000101111;
12'b010010111000: finv2 = 23'b00110001010101101110001;
12'b010010111001: finv2 = 23'b00110001001110010110101;
12'b010010111010: finv2 = 23'b00110001000110111111100;
12'b010010111011: finv2 = 23'b00110000111111101000100;
12'b010010111100: finv2 = 23'b00110000111000010001111;
12'b010010111101: finv2 = 23'b00110000110000111011100;
12'b010010111110: finv2 = 23'b00110000101001100101011;
12'b010010111111: finv2 = 23'b00110000100010001111100;
12'b010011000000: finv2 = 23'b00110000011010111001111;
12'b010011000001: finv2 = 23'b00110000010011100100100;
12'b010011000010: finv2 = 23'b00110000001100001111100;
12'b010011000011: finv2 = 23'b00110000000100111010101;
12'b010011000100: finv2 = 23'b00101111111101100110001;
12'b010011000101: finv2 = 23'b00101111110110010001111;
12'b010011000110: finv2 = 23'b00101111101110111101111;
12'b010011000111: finv2 = 23'b00101111100111101010001;
12'b010011001000: finv2 = 23'b00101111100000010110101;
12'b010011001001: finv2 = 23'b00101111011001000011011;
12'b010011001010: finv2 = 23'b00101111010001110000011;
12'b010011001011: finv2 = 23'b00101111001010011101110;
12'b010011001100: finv2 = 23'b00101111000011001011010;
12'b010011001101: finv2 = 23'b00101110111011111001001;
12'b010011001110: finv2 = 23'b00101110110100100111010;
12'b010011001111: finv2 = 23'b00101110101101010101101;
12'b010011010000: finv2 = 23'b00101110100110000100010;
12'b010011010001: finv2 = 23'b00101110011110110011001;
12'b010011010010: finv2 = 23'b00101110010111100010010;
12'b010011010011: finv2 = 23'b00101110010000010001101;
12'b010011010100: finv2 = 23'b00101110001001000001010;
12'b010011010101: finv2 = 23'b00101110000001110001010;
12'b010011010110: finv2 = 23'b00101101111010100001011;
12'b010011010111: finv2 = 23'b00101101110011010001111;
12'b010011011000: finv2 = 23'b00101101101100000010100;
12'b010011011001: finv2 = 23'b00101101100100110011100;
12'b010011011010: finv2 = 23'b00101101011101100100110;
12'b010011011011: finv2 = 23'b00101101010110010110010;
12'b010011011100: finv2 = 23'b00101101001111001000000;
12'b010011011101: finv2 = 23'b00101101000111111010000;
12'b010011011110: finv2 = 23'b00101101000000101100010;
12'b010011011111: finv2 = 23'b00101100111001011110110;
12'b010011100000: finv2 = 23'b00101100110010010001101;
12'b010011100001: finv2 = 23'b00101100101011000100101;
12'b010011100010: finv2 = 23'b00101100100011110111111;
12'b010011100011: finv2 = 23'b00101100011100101011100;
12'b010011100100: finv2 = 23'b00101100010101011111011;
12'b010011100101: finv2 = 23'b00101100001110010011011;
12'b010011100110: finv2 = 23'b00101100000111000111110;
12'b010011100111: finv2 = 23'b00101011111111111100011;
12'b010011101000: finv2 = 23'b00101011111000110001001;
12'b010011101001: finv2 = 23'b00101011110001100110010;
12'b010011101010: finv2 = 23'b00101011101010011011101;
12'b010011101011: finv2 = 23'b00101011100011010001010;
12'b010011101100: finv2 = 23'b00101011011100000111001;
12'b010011101101: finv2 = 23'b00101011010100111101010;
12'b010011101110: finv2 = 23'b00101011001101110011101;
12'b010011101111: finv2 = 23'b00101011000110101010011;
12'b010011110000: finv2 = 23'b00101010111111100001010;
12'b010011110001: finv2 = 23'b00101010111000011000011;
12'b010011110010: finv2 = 23'b00101010110001001111110;
12'b010011110011: finv2 = 23'b00101010101010000111100;
12'b010011110100: finv2 = 23'b00101010100010111111011;
12'b010011110101: finv2 = 23'b00101010011011110111101;
12'b010011110110: finv2 = 23'b00101010010100110000000;
12'b010011110111: finv2 = 23'b00101010001101101000110;
12'b010011111000: finv2 = 23'b00101010000110100001101;
12'b010011111001: finv2 = 23'b00101001111111011010111;
12'b010011111010: finv2 = 23'b00101001111000010100010;
12'b010011111011: finv2 = 23'b00101001110001001110000;
12'b010011111100: finv2 = 23'b00101001101010001000000;
12'b010011111101: finv2 = 23'b00101001100011000010010;
12'b010011111110: finv2 = 23'b00101001011011111100101;
12'b010011111111: finv2 = 23'b00101001010100110111011;
12'b010100000000: finv2 = 23'b00101001001101110010011;
12'b010100000001: finv2 = 23'b00101001000110101101101;
12'b010100000010: finv2 = 23'b00101000111111101001001;
12'b010100000011: finv2 = 23'b00101000111000100100110;
12'b010100000100: finv2 = 23'b00101000110001100000110;
12'b010100000101: finv2 = 23'b00101000101010011101000;
12'b010100000110: finv2 = 23'b00101000100011011001100;
12'b010100000111: finv2 = 23'b00101000011100010110010;
12'b010100001000: finv2 = 23'b00101000010101010011010;
12'b010100001001: finv2 = 23'b00101000001110010000100;
12'b010100001010: finv2 = 23'b00101000000111001110000;
12'b010100001011: finv2 = 23'b00101000000000001011110;
12'b010100001100: finv2 = 23'b00100111111001001001110;
12'b010100001101: finv2 = 23'b00100111110010001000000;
12'b010100001110: finv2 = 23'b00100111101011000110100;
12'b010100001111: finv2 = 23'b00100111100100000101010;
12'b010100010000: finv2 = 23'b00100111011101000100001;
12'b010100010001: finv2 = 23'b00100111010110000011011;
12'b010100010010: finv2 = 23'b00100111001111000010111;
12'b010100010011: finv2 = 23'b00100111001000000010101;
12'b010100010100: finv2 = 23'b00100111000001000010101;
12'b010100010101: finv2 = 23'b00100110111010000010111;
12'b010100010110: finv2 = 23'b00100110110011000011011;
12'b010100010111: finv2 = 23'b00100110101100000100001;
12'b010100011000: finv2 = 23'b00100110100101000101001;
12'b010100011001: finv2 = 23'b00100110011110000110011;
12'b010100011010: finv2 = 23'b00100110010111000111111;
12'b010100011011: finv2 = 23'b00100110010000001001101;
12'b010100011100: finv2 = 23'b00100110001001001011100;
12'b010100011101: finv2 = 23'b00100110000010001101110;
12'b010100011110: finv2 = 23'b00100101111011010000010;
12'b010100011111: finv2 = 23'b00100101110100010011000;
12'b010100100000: finv2 = 23'b00100101101101010110000;
12'b010100100001: finv2 = 23'b00100101100110011001001;
12'b010100100010: finv2 = 23'b00100101011111011100101;
12'b010100100011: finv2 = 23'b00100101011000100000011;
12'b010100100100: finv2 = 23'b00100101010001100100010;
12'b010100100101: finv2 = 23'b00100101001010101000100;
12'b010100100110: finv2 = 23'b00100101000011101101000;
12'b010100100111: finv2 = 23'b00100100111100110001101;
12'b010100101000: finv2 = 23'b00100100110101110110101;
12'b010100101001: finv2 = 23'b00100100101110111011110;
12'b010100101010: finv2 = 23'b00100100101000000001001;
12'b010100101011: finv2 = 23'b00100100100001000110111;
12'b010100101100: finv2 = 23'b00100100011010001100110;
12'b010100101101: finv2 = 23'b00100100010011010011000;
12'b010100101110: finv2 = 23'b00100100001100011001011;
12'b010100101111: finv2 = 23'b00100100000101100000000;
12'b010100110000: finv2 = 23'b00100011111110100110111;
12'b010100110001: finv2 = 23'b00100011110111101110000;
12'b010100110010: finv2 = 23'b00100011110000110101011;
12'b010100110011: finv2 = 23'b00100011101001111101000;
12'b010100110100: finv2 = 23'b00100011100011000100111;
12'b010100110101: finv2 = 23'b00100011011100001101000;
12'b010100110110: finv2 = 23'b00100011010101010101011;
12'b010100110111: finv2 = 23'b00100011001110011110000;
12'b010100111000: finv2 = 23'b00100011000111100110111;
12'b010100111001: finv2 = 23'b00100011000000101111111;
12'b010100111010: finv2 = 23'b00100010111001111001010;
12'b010100111011: finv2 = 23'b00100010110011000010110;
12'b010100111100: finv2 = 23'b00100010101100001100101;
12'b010100111101: finv2 = 23'b00100010100101010110101;
12'b010100111110: finv2 = 23'b00100010011110100001000;
12'b010100111111: finv2 = 23'b00100010010111101011100;
12'b010101000000: finv2 = 23'b00100010010000110110010;
12'b010101000001: finv2 = 23'b00100010001010000001010;
12'b010101000010: finv2 = 23'b00100010000011001100100;
12'b010101000011: finv2 = 23'b00100001111100011000000;
12'b010101000100: finv2 = 23'b00100001110101100011110;
12'b010101000101: finv2 = 23'b00100001101110101111110;
12'b010101000110: finv2 = 23'b00100001100111111100000;
12'b010101000111: finv2 = 23'b00100001100001001000100;
12'b010101001000: finv2 = 23'b00100001011010010101001;
12'b010101001001: finv2 = 23'b00100001010011100010001;
12'b010101001010: finv2 = 23'b00100001001100101111010;
12'b010101001011: finv2 = 23'b00100001000101111100110;
12'b010101001100: finv2 = 23'b00100000111111001010011;
12'b010101001101: finv2 = 23'b00100000111000011000010;
12'b010101001110: finv2 = 23'b00100000110001100110011;
12'b010101001111: finv2 = 23'b00100000101010110100110;
12'b010101010000: finv2 = 23'b00100000100100000011011;
12'b010101010001: finv2 = 23'b00100000011101010010010;
12'b010101010010: finv2 = 23'b00100000010110100001011;
12'b010101010011: finv2 = 23'b00100000001111110000101;
12'b010101010100: finv2 = 23'b00100000001001000000010;
12'b010101010101: finv2 = 23'b00100000000010010000000;
12'b010101010110: finv2 = 23'b00011111111011100000000;
12'b010101010111: finv2 = 23'b00011111110100110000011;
12'b010101011000: finv2 = 23'b00011111101110000000111;
12'b010101011001: finv2 = 23'b00011111100111010001101;
12'b010101011010: finv2 = 23'b00011111100000100010101;
12'b010101011011: finv2 = 23'b00011111011001110011110;
12'b010101011100: finv2 = 23'b00011111010011000101010;
12'b010101011101: finv2 = 23'b00011111001100010111000;
12'b010101011110: finv2 = 23'b00011111000101101000111;
12'b010101011111: finv2 = 23'b00011110111110111011000;
12'b010101100000: finv2 = 23'b00011110111000001101100;
12'b010101100001: finv2 = 23'b00011110110001100000001;
12'b010101100010: finv2 = 23'b00011110101010110011000;
12'b010101100011: finv2 = 23'b00011110100100000110001;
12'b010101100100: finv2 = 23'b00011110011101011001011;
12'b010101100101: finv2 = 23'b00011110010110101101000;
12'b010101100110: finv2 = 23'b00011110010000000000111;
12'b010101100111: finv2 = 23'b00011110001001010100111;
12'b010101101000: finv2 = 23'b00011110000010101001001;
12'b010101101001: finv2 = 23'b00011101111011111101101;
12'b010101101010: finv2 = 23'b00011101110101010010011;
12'b010101101011: finv2 = 23'b00011101101110100111011;
12'b010101101100: finv2 = 23'b00011101100111111100101;
12'b010101101101: finv2 = 23'b00011101100001010010001;
12'b010101101110: finv2 = 23'b00011101011010100111110;
12'b010101101111: finv2 = 23'b00011101010011111101101;
12'b010101110000: finv2 = 23'b00011101001101010011111;
12'b010101110001: finv2 = 23'b00011101000110101010010;
12'b010101110010: finv2 = 23'b00011101000000000000111;
12'b010101110011: finv2 = 23'b00011100111001010111101;
12'b010101110100: finv2 = 23'b00011100110010101110110;
12'b010101110101: finv2 = 23'b00011100101100000110001;
12'b010101110110: finv2 = 23'b00011100100101011101101;
12'b010101110111: finv2 = 23'b00011100011110110101011;
12'b010101111000: finv2 = 23'b00011100011000001101011;
12'b010101111001: finv2 = 23'b00011100010001100101101;
12'b010101111010: finv2 = 23'b00011100001010111110001;
12'b010101111011: finv2 = 23'b00011100000100010110110;
12'b010101111100: finv2 = 23'b00011011111101101111110;
12'b010101111101: finv2 = 23'b00011011110111001000111;
12'b010101111110: finv2 = 23'b00011011110000100010010;
12'b010101111111: finv2 = 23'b00011011101001111011111;
12'b010110000000: finv2 = 23'b00011011100011010101110;
12'b010110000001: finv2 = 23'b00011011011100101111111;
12'b010110000010: finv2 = 23'b00011011010110001010001;
12'b010110000011: finv2 = 23'b00011011001111100100110;
12'b010110000100: finv2 = 23'b00011011001000111111100;
12'b010110000101: finv2 = 23'b00011011000010011010100;
12'b010110000110: finv2 = 23'b00011010111011110101110;
12'b010110000111: finv2 = 23'b00011010110101010001001;
12'b010110001000: finv2 = 23'b00011010101110101100111;
12'b010110001001: finv2 = 23'b00011010101000001000110;
12'b010110001010: finv2 = 23'b00011010100001100100111;
12'b010110001011: finv2 = 23'b00011010011011000001010;
12'b010110001100: finv2 = 23'b00011010010100011101111;
12'b010110001101: finv2 = 23'b00011010001101111010110;
12'b010110001110: finv2 = 23'b00011010000111010111110;
12'b010110001111: finv2 = 23'b00011010000000110101001;
12'b010110010000: finv2 = 23'b00011001111010010010101;
12'b010110010001: finv2 = 23'b00011001110011110000011;
12'b010110010010: finv2 = 23'b00011001101101001110011;
12'b010110010011: finv2 = 23'b00011001100110101100100;
12'b010110010100: finv2 = 23'b00011001100000001010111;
12'b010110010101: finv2 = 23'b00011001011001101001101;
12'b010110010110: finv2 = 23'b00011001010011001000100;
12'b010110010111: finv2 = 23'b00011001001100100111100;
12'b010110011000: finv2 = 23'b00011001000110000110111;
12'b010110011001: finv2 = 23'b00011000111111100110100;
12'b010110011010: finv2 = 23'b00011000111001000110010;
12'b010110011011: finv2 = 23'b00011000110010100110010;
12'b010110011100: finv2 = 23'b00011000101100000110100;
12'b010110011101: finv2 = 23'b00011000100101100110111;
12'b010110011110: finv2 = 23'b00011000011111000111101;
12'b010110011111: finv2 = 23'b00011000011000101000100;
12'b010110100000: finv2 = 23'b00011000010010001001101;
12'b010110100001: finv2 = 23'b00011000001011101011000;
12'b010110100010: finv2 = 23'b00011000000101001100101;
12'b010110100011: finv2 = 23'b00010111111110101110011;
12'b010110100100: finv2 = 23'b00010111111000010000011;
12'b010110100101: finv2 = 23'b00010111110001110010101;
12'b010110100110: finv2 = 23'b00010111101011010101001;
12'b010110100111: finv2 = 23'b00010111100100110111111;
12'b010110101000: finv2 = 23'b00010111011110011010110;
12'b010110101001: finv2 = 23'b00010111010111111101111;
12'b010110101010: finv2 = 23'b00010111010001100001010;
12'b010110101011: finv2 = 23'b00010111001011000100111;
12'b010110101100: finv2 = 23'b00010111000100101000110;
12'b010110101101: finv2 = 23'b00010110111110001100110;
12'b010110101110: finv2 = 23'b00010110110111110001000;
12'b010110101111: finv2 = 23'b00010110110001010101100;
12'b010110110000: finv2 = 23'b00010110101010111010010;
12'b010110110001: finv2 = 23'b00010110100100011111001;
12'b010110110010: finv2 = 23'b00010110011110000100010;
12'b010110110011: finv2 = 23'b00010110010111101001101;
12'b010110110100: finv2 = 23'b00010110010001001111010;
12'b010110110101: finv2 = 23'b00010110001010110101001;
12'b010110110110: finv2 = 23'b00010110000100011011001;
12'b010110110111: finv2 = 23'b00010101111110000001011;
12'b010110111000: finv2 = 23'b00010101110111100111111;
12'b010110111001: finv2 = 23'b00010101110001001110101;
12'b010110111010: finv2 = 23'b00010101101010110101100;
12'b010110111011: finv2 = 23'b00010101100100011100101;
12'b010110111100: finv2 = 23'b00010101011110000100000;
12'b010110111101: finv2 = 23'b00010101010111101011101;
12'b010110111110: finv2 = 23'b00010101010001010011011;
12'b010110111111: finv2 = 23'b00010101001010111011011;
12'b010111000000: finv2 = 23'b00010101000100100011101;
12'b010111000001: finv2 = 23'b00010100111110001100001;
12'b010111000010: finv2 = 23'b00010100110111110100111;
12'b010111000011: finv2 = 23'b00010100110001011101110;
12'b010111000100: finv2 = 23'b00010100101011000110111;
12'b010111000101: finv2 = 23'b00010100100100110000010;
12'b010111000110: finv2 = 23'b00010100011110011001110;
12'b010111000111: finv2 = 23'b00010100011000000011100;
12'b010111001000: finv2 = 23'b00010100010001101101100;
12'b010111001001: finv2 = 23'b00010100001011010111110;
12'b010111001010: finv2 = 23'b00010100000101000010010;
12'b010111001011: finv2 = 23'b00010011111110101100111;
12'b010111001100: finv2 = 23'b00010011111000010111110;
12'b010111001101: finv2 = 23'b00010011110010000010110;
12'b010111001110: finv2 = 23'b00010011101011101110001;
12'b010111001111: finv2 = 23'b00010011100101011001101;
12'b010111010000: finv2 = 23'b00010011011111000101011;
12'b010111010001: finv2 = 23'b00010011011000110001011;
12'b010111010010: finv2 = 23'b00010011010010011101100;
12'b010111010011: finv2 = 23'b00010011001100001001111;
12'b010111010100: finv2 = 23'b00010011000101110110100;
12'b010111010101: finv2 = 23'b00010010111111100011011;
12'b010111010110: finv2 = 23'b00010010111001010000011;
12'b010111010111: finv2 = 23'b00010010110010111101101;
12'b010111011000: finv2 = 23'b00010010101100101011001;
12'b010111011001: finv2 = 23'b00010010100110011000110;
12'b010111011010: finv2 = 23'b00010010100000000110110;
12'b010111011011: finv2 = 23'b00010010011001110100110;
12'b010111011100: finv2 = 23'b00010010010011100011001;
12'b010111011101: finv2 = 23'b00010010001101010001110;
12'b010111011110: finv2 = 23'b00010010000111000000100;
12'b010111011111: finv2 = 23'b00010010000000101111100;
12'b010111100000: finv2 = 23'b00010001111010011110101;
12'b010111100001: finv2 = 23'b00010001110100001110000;
12'b010111100010: finv2 = 23'b00010001101101111101101;
12'b010111100011: finv2 = 23'b00010001100111101101100;
12'b010111100100: finv2 = 23'b00010001100001011101101;
12'b010111100101: finv2 = 23'b00010001011011001101111;
12'b010111100110: finv2 = 23'b00010001010100111110011;
12'b010111100111: finv2 = 23'b00010001001110101111000;
12'b010111101000: finv2 = 23'b00010001001000011111111;
12'b010111101001: finv2 = 23'b00010001000010010001000;
12'b010111101010: finv2 = 23'b00010000111100000010011;
12'b010111101011: finv2 = 23'b00010000110101110011111;
12'b010111101100: finv2 = 23'b00010000101111100101110;
12'b010111101101: finv2 = 23'b00010000101001010111101;
12'b010111101110: finv2 = 23'b00010000100011001001111;
12'b010111101111: finv2 = 23'b00010000011100111100010;
12'b010111110000: finv2 = 23'b00010000010110101110111;
12'b010111110001: finv2 = 23'b00010000010000100001110;
12'b010111110010: finv2 = 23'b00010000001010010100110;
12'b010111110011: finv2 = 23'b00010000000100001000000;
12'b010111110100: finv2 = 23'b00001111111101111011011;
12'b010111110101: finv2 = 23'b00001111110111101111001;
12'b010111110110: finv2 = 23'b00001111110001100011000;
12'b010111110111: finv2 = 23'b00001111101011010111001;
12'b010111111000: finv2 = 23'b00001111100101001011011;
12'b010111111001: finv2 = 23'b00001111011110111111111;
12'b010111111010: finv2 = 23'b00001111011000110100101;
12'b010111111011: finv2 = 23'b00001111010010101001101;
12'b010111111100: finv2 = 23'b00001111001100011110110;
12'b010111111101: finv2 = 23'b00001111000110010100001;
12'b010111111110: finv2 = 23'b00001111000000001001101;
12'b010111111111: finv2 = 23'b00001110111001111111011;
12'b011000000000: finv2 = 23'b00001110110011110101011;
12'b011000000001: finv2 = 23'b00001110101101101011101;
12'b011000000010: finv2 = 23'b00001110100111100010000;
12'b011000000011: finv2 = 23'b00001110100001011000101;
12'b011000000100: finv2 = 23'b00001110011011001111100;
12'b011000000101: finv2 = 23'b00001110010101000110100;
12'b011000000110: finv2 = 23'b00001110001110111101110;
12'b011000000111: finv2 = 23'b00001110001000110101010;
12'b011000001000: finv2 = 23'b00001110000010101100111;
12'b011000001001: finv2 = 23'b00001101111100100100110;
12'b011000001010: finv2 = 23'b00001101110110011100111;
12'b011000001011: finv2 = 23'b00001101110000010101001;
12'b011000001100: finv2 = 23'b00001101101010001101101;
12'b011000001101: finv2 = 23'b00001101100100000110011;
12'b011000001110: finv2 = 23'b00001101011101111111010;
12'b011000001111: finv2 = 23'b00001101010111111000011;
12'b011000010000: finv2 = 23'b00001101010001110001110;
12'b011000010001: finv2 = 23'b00001101001011101011010;
12'b011000010010: finv2 = 23'b00001101000101100101000;
12'b011000010011: finv2 = 23'b00001100111111011110111;
12'b011000010100: finv2 = 23'b00001100111001011001001;
12'b011000010101: finv2 = 23'b00001100110011010011100;
12'b011000010110: finv2 = 23'b00001100101101001110000;
12'b011000010111: finv2 = 23'b00001100100111001000110;
12'b011000011000: finv2 = 23'b00001100100001000011110;
12'b011000011001: finv2 = 23'b00001100011010111111000;
12'b011000011010: finv2 = 23'b00001100010100111010011;
12'b011000011011: finv2 = 23'b00001100001110110110000;
12'b011000011100: finv2 = 23'b00001100001000110001110;
12'b011000011101: finv2 = 23'b00001100000010101101110;
12'b011000011110: finv2 = 23'b00001011111100101010000;
12'b011000011111: finv2 = 23'b00001011110110100110100;
12'b011000100000: finv2 = 23'b00001011110000100011001;
12'b011000100001: finv2 = 23'b00001011101010011111111;
12'b011000100010: finv2 = 23'b00001011100100011101000;
12'b011000100011: finv2 = 23'b00001011011110011010010;
12'b011000100100: finv2 = 23'b00001011011000010111101;
12'b011000100101: finv2 = 23'b00001011010010010101010;
12'b011000100110: finv2 = 23'b00001011001100010011001;
12'b011000100111: finv2 = 23'b00001011000110010001010;
12'b011000101000: finv2 = 23'b00001011000000001111100;
12'b011000101001: finv2 = 23'b00001010111010001110000;
12'b011000101010: finv2 = 23'b00001010110100001100101;
12'b011000101011: finv2 = 23'b00001010101110001011100;
12'b011000101100: finv2 = 23'b00001010101000001010101;
12'b011000101101: finv2 = 23'b00001010100010001001111;
12'b011000101110: finv2 = 23'b00001010011100001001011;
12'b011000101111: finv2 = 23'b00001010010110001001001;
12'b011000110000: finv2 = 23'b00001010010000001001000;
12'b011000110001: finv2 = 23'b00001010001010001001000;
12'b011000110010: finv2 = 23'b00001010000100001001011;
12'b011000110011: finv2 = 23'b00001001111110001001111;
12'b011000110100: finv2 = 23'b00001001111000001010101;
12'b011000110101: finv2 = 23'b00001001110010001011100;
12'b011000110110: finv2 = 23'b00001001101100001100101;
12'b011000110111: finv2 = 23'b00001001100110001101111;
12'b011000111000: finv2 = 23'b00001001100000001111011;
12'b011000111001: finv2 = 23'b00001001011010010001001;
12'b011000111010: finv2 = 23'b00001001010100010011000;
12'b011000111011: finv2 = 23'b00001001001110010101001;
12'b011000111100: finv2 = 23'b00001001001000010111100;
12'b011000111101: finv2 = 23'b00001001000010011010000;
12'b011000111110: finv2 = 23'b00001000111100011100110;
12'b011000111111: finv2 = 23'b00001000110110011111101;
12'b011001000000: finv2 = 23'b00001000110000100010110;
12'b011001000001: finv2 = 23'b00001000101010100110001;
12'b011001000010: finv2 = 23'b00001000100100101001101;
12'b011001000011: finv2 = 23'b00001000011110101101011;
12'b011001000100: finv2 = 23'b00001000011000110001010;
12'b011001000101: finv2 = 23'b00001000010010110101011;
12'b011001000110: finv2 = 23'b00001000001100111001110;
12'b011001000111: finv2 = 23'b00001000000110111110010;
12'b011001001000: finv2 = 23'b00001000000001000011000;
12'b011001001001: finv2 = 23'b00000111111011000111111;
12'b011001001010: finv2 = 23'b00000111110101001101000;
12'b011001001011: finv2 = 23'b00000111101111010010011;
12'b011001001100: finv2 = 23'b00000111101001010111111;
12'b011001001101: finv2 = 23'b00000111100011011101101;
12'b011001001110: finv2 = 23'b00000111011101100011100;
12'b011001001111: finv2 = 23'b00000111010111101001101;
12'b011001010000: finv2 = 23'b00000111010001101111111;
12'b011001010001: finv2 = 23'b00000111001011110110100;
12'b011001010010: finv2 = 23'b00000111000101111101001;
12'b011001010011: finv2 = 23'b00000111000000000100001;
12'b011001010100: finv2 = 23'b00000110111010001011001;
12'b011001010101: finv2 = 23'b00000110110100010010100;
12'b011001010110: finv2 = 23'b00000110101110011010000;
12'b011001010111: finv2 = 23'b00000110101000100001101;
12'b011001011000: finv2 = 23'b00000110100010101001101;
12'b011001011001: finv2 = 23'b00000110011100110001101;
12'b011001011010: finv2 = 23'b00000110010110111010000;
12'b011001011011: finv2 = 23'b00000110010001000010100;
12'b011001011100: finv2 = 23'b00000110001011001011001;
12'b011001011101: finv2 = 23'b00000110000101010100000;
12'b011001011110: finv2 = 23'b00000101111111011101001;
12'b011001011111: finv2 = 23'b00000101111001100110011;
12'b011001100000: finv2 = 23'b00000101110011101111111;
12'b011001100001: finv2 = 23'b00000101101101111001100;
12'b011001100010: finv2 = 23'b00000101101000000011011;
12'b011001100011: finv2 = 23'b00000101100010001101100;
12'b011001100100: finv2 = 23'b00000101011100010111110;
12'b011001100101: finv2 = 23'b00000101010110100010001;
12'b011001100110: finv2 = 23'b00000101010000101100110;
12'b011001100111: finv2 = 23'b00000101001010110111101;
12'b011001101000: finv2 = 23'b00000101000101000010101;
12'b011001101001: finv2 = 23'b00000100111111001101111;
12'b011001101010: finv2 = 23'b00000100111001011001011;
12'b011001101011: finv2 = 23'b00000100110011100101000;
12'b011001101100: finv2 = 23'b00000100101101110000110;
12'b011001101101: finv2 = 23'b00000100100111111100110;
12'b011001101110: finv2 = 23'b00000100100010001001000;
12'b011001101111: finv2 = 23'b00000100011100010101011;
12'b011001110000: finv2 = 23'b00000100010110100010000;
12'b011001110001: finv2 = 23'b00000100010000101110110;
12'b011001110010: finv2 = 23'b00000100001010111011110;
12'b011001110011: finv2 = 23'b00000100000101001000111;
12'b011001110100: finv2 = 23'b00000011111111010110010;
12'b011001110101: finv2 = 23'b00000011111001100011111;
12'b011001110110: finv2 = 23'b00000011110011110001101;
12'b011001110111: finv2 = 23'b00000011101101111111100;
12'b011001111000: finv2 = 23'b00000011101000001101110;
12'b011001111001: finv2 = 23'b00000011100010011100000;
12'b011001111010: finv2 = 23'b00000011011100101010100;
12'b011001111011: finv2 = 23'b00000011010110111001010;
12'b011001111100: finv2 = 23'b00000011010001001000001;
12'b011001111101: finv2 = 23'b00000011001011010111010;
12'b011001111110: finv2 = 23'b00000011000101100110101;
12'b011001111111: finv2 = 23'b00000010111111110110001;
12'b011010000000: finv2 = 23'b00000010111010000101110;
12'b011010000001: finv2 = 23'b00000010110100010101101;
12'b011010000010: finv2 = 23'b00000010101110100101101;
12'b011010000011: finv2 = 23'b00000010101000110110000;
12'b011010000100: finv2 = 23'b00000010100011000110011;
12'b011010000101: finv2 = 23'b00000010011101010111000;
12'b011010000110: finv2 = 23'b00000010010111100111111;
12'b011010000111: finv2 = 23'b00000010010001111000111;
12'b011010001000: finv2 = 23'b00000010001100001010001;
12'b011010001001: finv2 = 23'b00000010000110011011100;
12'b011010001010: finv2 = 23'b00000010000000101101001;
12'b011010001011: finv2 = 23'b00000001111010111110111;
12'b011010001100: finv2 = 23'b00000001110101010000111;
12'b011010001101: finv2 = 23'b00000001101111100011000;
12'b011010001110: finv2 = 23'b00000001101001110101011;
12'b011010001111: finv2 = 23'b00000001100100000111111;
12'b011010010000: finv2 = 23'b00000001011110011010101;
12'b011010010001: finv2 = 23'b00000001011000101101100;
12'b011010010010: finv2 = 23'b00000001010011000000101;
12'b011010010011: finv2 = 23'b00000001001101010100000;
12'b011010010100: finv2 = 23'b00000001000111100111100;
12'b011010010101: finv2 = 23'b00000001000001111011001;
12'b011010010110: finv2 = 23'b00000000111100001111000;
12'b011010010111: finv2 = 23'b00000000110110100011000;
12'b011010011000: finv2 = 23'b00000000110000110111010;
12'b011010011001: finv2 = 23'b00000000101011001011110;
12'b011010011010: finv2 = 23'b00000000100101100000011;
12'b011010011011: finv2 = 23'b00000000011111110101001;
12'b011010011100: finv2 = 23'b00000000011010001010001;
12'b011010011101: finv2 = 23'b00000000010100011111011;
12'b011010011110: finv2 = 23'b00000000001110110100110;
12'b011010011111: finv2 = 23'b00000000001001001010010;
12'b011010100000: finv2 = 23'b00000000000011100000000;
12'b011010100001: finv2 = 23'b11111111111011101100000;
12'b011010100010: finv2 = 23'b11111111110000011000010;
12'b011010100011: finv2 = 23'b11111111100101000100111;
12'b011010100100: finv2 = 23'b11111111011001110001111;
12'b011010100101: finv2 = 23'b11111111001110011111010;
12'b011010100110: finv2 = 23'b11111111000011001101000;
12'b011010100111: finv2 = 23'b11111110110111111011001;
12'b011010101000: finv2 = 23'b11111110101100101001101;
12'b011010101001: finv2 = 23'b11111110100001011000100;
12'b011010101010: finv2 = 23'b11111110010110000111110;
12'b011010101011: finv2 = 23'b11111110001010110111011;
12'b011010101100: finv2 = 23'b11111101111111100111011;
12'b011010101101: finv2 = 23'b11111101110100010111101;
12'b011010101110: finv2 = 23'b11111101101001001000011;
12'b011010101111: finv2 = 23'b11111101011101111001100;
12'b011010110000: finv2 = 23'b11111101010010101011000;
12'b011010110001: finv2 = 23'b11111101000111011100111;
12'b011010110010: finv2 = 23'b11111100111100001111000;
12'b011010110011: finv2 = 23'b11111100110001000001101;
12'b011010110100: finv2 = 23'b11111100100101110100101;
12'b011010110101: finv2 = 23'b11111100011010100111111;
12'b011010110110: finv2 = 23'b11111100001111011011101;
12'b011010110111: finv2 = 23'b11111100000100001111101;
12'b011010111000: finv2 = 23'b11111011111001000100001;
12'b011010111001: finv2 = 23'b11111011101101111000111;
12'b011010111010: finv2 = 23'b11111011100010101110001;
12'b011010111011: finv2 = 23'b11111011010111100011101;
12'b011010111100: finv2 = 23'b11111011001100011001100;
12'b011010111101: finv2 = 23'b11111011000001001111111;
12'b011010111110: finv2 = 23'b11111010110110000110100;
12'b011010111111: finv2 = 23'b11111010101010111101100;
12'b011011000000: finv2 = 23'b11111010011111110100111;
12'b011011000001: finv2 = 23'b11111010010100101100101;
12'b011011000010: finv2 = 23'b11111010001001100100110;
12'b011011000011: finv2 = 23'b11111001111110011101010;
12'b011011000100: finv2 = 23'b11111001110011010110000;
12'b011011000101: finv2 = 23'b11111001101000001111010;
12'b011011000110: finv2 = 23'b11111001011101001000111;
12'b011011000111: finv2 = 23'b11111001010010000010110;
12'b011011001000: finv2 = 23'b11111001000110111101001;
12'b011011001001: finv2 = 23'b11111000111011110111110;
12'b011011001010: finv2 = 23'b11111000110000110010111;
12'b011011001011: finv2 = 23'b11111000100101101110010;
12'b011011001100: finv2 = 23'b11111000011010101010000;
12'b011011001101: finv2 = 23'b11111000001111100110001;
12'b011011001110: finv2 = 23'b11111000000100100010101;
12'b011011001111: finv2 = 23'b11110111111001011111100;
12'b011011010000: finv2 = 23'b11110111101110011100110;
12'b011011010001: finv2 = 23'b11110111100011011010010;
12'b011011010010: finv2 = 23'b11110111011000011000010;
12'b011011010011: finv2 = 23'b11110111001101010110100;
12'b011011010100: finv2 = 23'b11110111000010010101010;
12'b011011010101: finv2 = 23'b11110110110111010100010;
12'b011011010110: finv2 = 23'b11110110101100010011101;
12'b011011010111: finv2 = 23'b11110110100001010011011;
12'b011011011000: finv2 = 23'b11110110010110010011100;
12'b011011011001: finv2 = 23'b11110110001011010100000;
12'b011011011010: finv2 = 23'b11110110000000010100111;
12'b011011011011: finv2 = 23'b11110101110101010110000;
12'b011011011100: finv2 = 23'b11110101101010010111101;
12'b011011011101: finv2 = 23'b11110101011111011001100;
12'b011011011110: finv2 = 23'b11110101010100011011111;
12'b011011011111: finv2 = 23'b11110101001001011110100;
12'b011011100000: finv2 = 23'b11110100111110100001100;
12'b011011100001: finv2 = 23'b11110100110011100100111;
12'b011011100010: finv2 = 23'b11110100101000101000100;
12'b011011100011: finv2 = 23'b11110100011101101100101;
12'b011011100100: finv2 = 23'b11110100010010110001000;
12'b011011100101: finv2 = 23'b11110100000111110101111;
12'b011011100110: finv2 = 23'b11110011111100111011000;
12'b011011100111: finv2 = 23'b11110011110010000000100;
12'b011011101000: finv2 = 23'b11110011100111000110011;
12'b011011101001: finv2 = 23'b11110011011100001100101;
12'b011011101010: finv2 = 23'b11110011010001010011001;
12'b011011101011: finv2 = 23'b11110011000110011010001;
12'b011011101100: finv2 = 23'b11110010111011100001011;
12'b011011101101: finv2 = 23'b11110010110000101001000;
12'b011011101110: finv2 = 23'b11110010100101110001000;
12'b011011101111: finv2 = 23'b11110010011010111001011;
12'b011011110000: finv2 = 23'b11110010010000000010001;
12'b011011110001: finv2 = 23'b11110010000101001011010;
12'b011011110010: finv2 = 23'b11110001111010010100101;
12'b011011110011: finv2 = 23'b11110001101111011110011;
12'b011011110100: finv2 = 23'b11110001100100101000100;
12'b011011110101: finv2 = 23'b11110001011001110011000;
12'b011011110110: finv2 = 23'b11110001001110111101111;
12'b011011110111: finv2 = 23'b11110001000100001001000;
12'b011011111000: finv2 = 23'b11110000111001010100101;
12'b011011111001: finv2 = 23'b11110000101110100000100;
12'b011011111010: finv2 = 23'b11110000100011101100110;
12'b011011111011: finv2 = 23'b11110000011000111001011;
12'b011011111100: finv2 = 23'b11110000001110000110011;
12'b011011111101: finv2 = 23'b11110000000011010011101;
12'b011011111110: finv2 = 23'b11101111111000100001011;
12'b011011111111: finv2 = 23'b11101111101101101111011;
12'b011100000000: finv2 = 23'b11101111100010111101110;
12'b011100000001: finv2 = 23'b11101111011000001100011;
12'b011100000010: finv2 = 23'b11101111001101011011100;
12'b011100000011: finv2 = 23'b11101111000010101010111;
12'b011100000100: finv2 = 23'b11101110110111111010101;
12'b011100000101: finv2 = 23'b11101110101101001010110;
12'b011100000110: finv2 = 23'b11101110100010011011010;
12'b011100000111: finv2 = 23'b11101110010111101100001;
12'b011100001000: finv2 = 23'b11101110001100111101010;
12'b011100001001: finv2 = 23'b11101110000010001110110;
12'b011100001010: finv2 = 23'b11101101110111100000101;
12'b011100001011: finv2 = 23'b11101101101100110010111;
12'b011100001100: finv2 = 23'b11101101100010000101100;
12'b011100001101: finv2 = 23'b11101101010111011000011;
12'b011100001110: finv2 = 23'b11101101001100101011101;
12'b011100001111: finv2 = 23'b11101101000001111111010;
12'b011100010000: finv2 = 23'b11101100110111010011010;
12'b011100010001: finv2 = 23'b11101100101100100111100;
12'b011100010010: finv2 = 23'b11101100100001111100001;
12'b011100010011: finv2 = 23'b11101100010111010001001;
12'b011100010100: finv2 = 23'b11101100001100100110100;
12'b011100010101: finv2 = 23'b11101100000001111100010;
12'b011100010110: finv2 = 23'b11101011110111010010010;
12'b011100010111: finv2 = 23'b11101011101100101000101;
12'b011100011000: finv2 = 23'b11101011100001111111011;
12'b011100011001: finv2 = 23'b11101011010111010110100;
12'b011100011010: finv2 = 23'b11101011001100101101111;
12'b011100011011: finv2 = 23'b11101011000010000101101;
12'b011100011100: finv2 = 23'b11101010110111011101110;
12'b011100011101: finv2 = 23'b11101010101100110110010;
12'b011100011110: finv2 = 23'b11101010100010001111000;
12'b011100011111: finv2 = 23'b11101010010111101000010;
12'b011100100000: finv2 = 23'b11101010001101000001101;
12'b011100100001: finv2 = 23'b11101010000010011011100;
12'b011100100010: finv2 = 23'b11101001110111110101110;
12'b011100100011: finv2 = 23'b11101001101101010000010;
12'b011100100100: finv2 = 23'b11101001100010101011001;
12'b011100100101: finv2 = 23'b11101001011000000110010;
12'b011100100110: finv2 = 23'b11101001001101100001111;
12'b011100100111: finv2 = 23'b11101001000010111101110;
12'b011100101000: finv2 = 23'b11101000111000011010000;
12'b011100101001: finv2 = 23'b11101000101101110110100;
12'b011100101010: finv2 = 23'b11101000100011010011100;
12'b011100101011: finv2 = 23'b11101000011000110000110;
12'b011100101100: finv2 = 23'b11101000001110001110011;
12'b011100101101: finv2 = 23'b11101000000011101100010;
12'b011100101110: finv2 = 23'b11100111111001001010101;
12'b011100101111: finv2 = 23'b11100111101110101001001;
12'b011100110000: finv2 = 23'b11100111100100001000001;
12'b011100110001: finv2 = 23'b11100111011001100111100;
12'b011100110010: finv2 = 23'b11100111001111000111001;
12'b011100110011: finv2 = 23'b11100111000100100111001;
12'b011100110100: finv2 = 23'b11100110111010000111011;
12'b011100110101: finv2 = 23'b11100110101111101000001;
12'b011100110110: finv2 = 23'b11100110100101001001001;
12'b011100110111: finv2 = 23'b11100110011010101010011;
12'b011100111000: finv2 = 23'b11100110010000001100001;
12'b011100111001: finv2 = 23'b11100110000101101110001;
12'b011100111010: finv2 = 23'b11100101111011010000100;
12'b011100111011: finv2 = 23'b11100101110000110011001;
12'b011100111100: finv2 = 23'b11100101100110010110001;
12'b011100111101: finv2 = 23'b11100101011011111001100;
12'b011100111110: finv2 = 23'b11100101010001011101010;
12'b011100111111: finv2 = 23'b11100101000111000001010;
12'b011101000000: finv2 = 23'b11100100111100100101101;
12'b011101000001: finv2 = 23'b11100100110010001010011;
12'b011101000010: finv2 = 23'b11100100100111101111100;
12'b011101000011: finv2 = 23'b11100100011101010100111;
12'b011101000100: finv2 = 23'b11100100010010111010100;
12'b011101000101: finv2 = 23'b11100100001000100000101;
12'b011101000110: finv2 = 23'b11100011111110000111000;
12'b011101000111: finv2 = 23'b11100011110011101101110;
12'b011101001000: finv2 = 23'b11100011101001010100110;
12'b011101001001: finv2 = 23'b11100011011110111100010;
12'b011101001010: finv2 = 23'b11100011010100100011111;
12'b011101001011: finv2 = 23'b11100011001010001100000;
12'b011101001100: finv2 = 23'b11100010111111110100011;
12'b011101001101: finv2 = 23'b11100010110101011101001;
12'b011101001110: finv2 = 23'b11100010101011000110010;
12'b011101001111: finv2 = 23'b11100010100000101111101;
12'b011101010000: finv2 = 23'b11100010010110011001011;
12'b011101010001: finv2 = 23'b11100010001100000011011;
12'b011101010010: finv2 = 23'b11100010000001101101110;
12'b011101010011: finv2 = 23'b11100001110111011000100;
12'b011101010100: finv2 = 23'b11100001101101000011101;
12'b011101010101: finv2 = 23'b11100001100010101111000;
12'b011101010110: finv2 = 23'b11100001011000011010110;
12'b011101010111: finv2 = 23'b11100001001110000110110;
12'b011101011000: finv2 = 23'b11100001000011110011001;
12'b011101011001: finv2 = 23'b11100000111001011111111;
12'b011101011010: finv2 = 23'b11100000101111001101000;
12'b011101011011: finv2 = 23'b11100000100100111010011;
12'b011101011100: finv2 = 23'b11100000011010101000000;
12'b011101011101: finv2 = 23'b11100000010000010110001;
12'b011101011110: finv2 = 23'b11100000000110000100100;
12'b011101011111: finv2 = 23'b11011111111011110011001;
12'b011101100000: finv2 = 23'b11011111110001100010001;
12'b011101100001: finv2 = 23'b11011111100111010001100;
12'b011101100010: finv2 = 23'b11011111011101000001010;
12'b011101100011: finv2 = 23'b11011111010010110001010;
12'b011101100100: finv2 = 23'b11011111001000100001101;
12'b011101100101: finv2 = 23'b11011110111110010010010;
12'b011101100110: finv2 = 23'b11011110110100000011010;
12'b011101100111: finv2 = 23'b11011110101001110100101;
12'b011101101000: finv2 = 23'b11011110011111100110010;
12'b011101101001: finv2 = 23'b11011110010101011000010;
12'b011101101010: finv2 = 23'b11011110001011001010101;
12'b011101101011: finv2 = 23'b11011110000000111101010;
12'b011101101100: finv2 = 23'b11011101110110110000010;
12'b011101101101: finv2 = 23'b11011101101100100011100;
12'b011101101110: finv2 = 23'b11011101100010010111001;
12'b011101101111: finv2 = 23'b11011101011000001011001;
12'b011101110000: finv2 = 23'b11011101001101111111011;
12'b011101110001: finv2 = 23'b11011101000011110100000;
12'b011101110010: finv2 = 23'b11011100111001101000111;
12'b011101110011: finv2 = 23'b11011100101111011110001;
12'b011101110100: finv2 = 23'b11011100100101010011110;
12'b011101110101: finv2 = 23'b11011100011011001001101;
12'b011101110110: finv2 = 23'b11011100010000111111111;
12'b011101110111: finv2 = 23'b11011100000110110110011;
12'b011101111000: finv2 = 23'b11011011111100101101010;
12'b011101111001: finv2 = 23'b11011011110010100100100;
12'b011101111010: finv2 = 23'b11011011101000011100000;
12'b011101111011: finv2 = 23'b11011011011110010011111;
12'b011101111100: finv2 = 23'b11011011010100001100000;
12'b011101111101: finv2 = 23'b11011011001010000100100;
12'b011101111110: finv2 = 23'b11011010111111111101010;
12'b011101111111: finv2 = 23'b11011010110101110110011;
12'b011110000000: finv2 = 23'b11011010101011101111111;
12'b011110000001: finv2 = 23'b11011010100001101001101;
12'b011110000010: finv2 = 23'b11011010010111100011110;
12'b011110000011: finv2 = 23'b11011010001101011110010;
12'b011110000100: finv2 = 23'b11011010000011011001000;
12'b011110000101: finv2 = 23'b11011001111001010100000;
12'b011110000110: finv2 = 23'b11011001101111001111011;
12'b011110000111: finv2 = 23'b11011001100101001011001;
12'b011110001000: finv2 = 23'b11011001011011000111001;
12'b011110001001: finv2 = 23'b11011001010001000011100;
12'b011110001010: finv2 = 23'b11011001000111000000010;
12'b011110001011: finv2 = 23'b11011000111100111101010;
12'b011110001100: finv2 = 23'b11011000110010111010100;
12'b011110001101: finv2 = 23'b11011000101000111000001;
12'b011110001110: finv2 = 23'b11011000011110110110001;
12'b011110001111: finv2 = 23'b11011000010100110100011;
12'b011110010000: finv2 = 23'b11011000001010110011000;
12'b011110010001: finv2 = 23'b11011000000000110001111;
12'b011110010010: finv2 = 23'b11010111110110110001001;
12'b011110010011: finv2 = 23'b11010111101100110000101;
12'b011110010100: finv2 = 23'b11010111100010110000100;
12'b011110010101: finv2 = 23'b11010111011000110000110;
12'b011110010110: finv2 = 23'b11010111001110110001010;
12'b011110010111: finv2 = 23'b11010111000100110010000;
12'b011110011000: finv2 = 23'b11010110111010110011001;
12'b011110011001: finv2 = 23'b11010110110000110100101;
12'b011110011010: finv2 = 23'b11010110100110110110011;
12'b011110011011: finv2 = 23'b11010110011100111000100;
12'b011110011100: finv2 = 23'b11010110010010111010111;
12'b011110011101: finv2 = 23'b11010110001000111101101;
12'b011110011110: finv2 = 23'b11010101111111000000101;
12'b011110011111: finv2 = 23'b11010101110101000100000;
12'b011110100000: finv2 = 23'b11010101101011000111101;
12'b011110100001: finv2 = 23'b11010101100001001011101;
12'b011110100010: finv2 = 23'b11010101010111010000000;
12'b011110100011: finv2 = 23'b11010101001101010100101;
12'b011110100100: finv2 = 23'b11010101000011011001100;
12'b011110100101: finv2 = 23'b11010100111001011110110;
12'b011110100110: finv2 = 23'b11010100101111100100011;
12'b011110100111: finv2 = 23'b11010100100101101010010;
12'b011110101000: finv2 = 23'b11010100011011110000011;
12'b011110101001: finv2 = 23'b11010100010001110110111;
12'b011110101010: finv2 = 23'b11010100000111111101110;
12'b011110101011: finv2 = 23'b11010011111110000100111;
12'b011110101100: finv2 = 23'b11010011110100001100010;
12'b011110101101: finv2 = 23'b11010011101010010100000;
12'b011110101110: finv2 = 23'b11010011100000011100001;
12'b011110101111: finv2 = 23'b11010011010110100100100;
12'b011110110000: finv2 = 23'b11010011001100101101001;
12'b011110110001: finv2 = 23'b11010011000010110110001;
12'b011110110010: finv2 = 23'b11010010111000111111100;
12'b011110110011: finv2 = 23'b11010010101111001001001;
12'b011110110100: finv2 = 23'b11010010100101010011001;
12'b011110110101: finv2 = 23'b11010010011011011101011;
12'b011110110110: finv2 = 23'b11010010010001100111111;
12'b011110110111: finv2 = 23'b11010010000111110010110;
12'b011110111000: finv2 = 23'b11010001111101111110000;
12'b011110111001: finv2 = 23'b11010001110100001001100;
12'b011110111010: finv2 = 23'b11010001101010010101010;
12'b011110111011: finv2 = 23'b11010001100000100001011;
12'b011110111100: finv2 = 23'b11010001010110101101110;
12'b011110111101: finv2 = 23'b11010001001100111010100;
12'b011110111110: finv2 = 23'b11010001000011000111101;
12'b011110111111: finv2 = 23'b11010000111001010101000;
12'b011111000000: finv2 = 23'b11010000101111100010101;
12'b011111000001: finv2 = 23'b11010000100101110000101;
12'b011111000010: finv2 = 23'b11010000011011111110111;
12'b011111000011: finv2 = 23'b11010000010010001101100;
12'b011111000100: finv2 = 23'b11010000001000011100011;
12'b011111000101: finv2 = 23'b11001111111110101011101;
12'b011111000110: finv2 = 23'b11001111110100111011001;
12'b011111000111: finv2 = 23'b11001111101011001010111;
12'b011111001000: finv2 = 23'b11001111100001011011000;
12'b011111001001: finv2 = 23'b11001111010111101011100;
12'b011111001010: finv2 = 23'b11001111001101111100010;
12'b011111001011: finv2 = 23'b11001111000100001101010;
12'b011111001100: finv2 = 23'b11001110111010011110101;
12'b011111001101: finv2 = 23'b11001110110000110000010;
12'b011111001110: finv2 = 23'b11001110100111000010010;
12'b011111001111: finv2 = 23'b11001110011101010100100;
12'b011111010000: finv2 = 23'b11001110010011100111001;
12'b011111010001: finv2 = 23'b11001110001001111010000;
12'b011111010010: finv2 = 23'b11001110000000001101010;
12'b011111010011: finv2 = 23'b11001101110110100000110;
12'b011111010100: finv2 = 23'b11001101101100110100100;
12'b011111010101: finv2 = 23'b11001101100011001000101;
12'b011111010110: finv2 = 23'b11001101011001011101001;
12'b011111010111: finv2 = 23'b11001101001111110001110;
12'b011111011000: finv2 = 23'b11001101000110000110111;
12'b011111011001: finv2 = 23'b11001100111100011100001;
12'b011111011010: finv2 = 23'b11001100110010110001110;
12'b011111011011: finv2 = 23'b11001100101001000111110;
12'b011111011100: finv2 = 23'b11001100011111011110000;
12'b011111011101: finv2 = 23'b11001100010101110100100;
12'b011111011110: finv2 = 23'b11001100001100001011011;
12'b011111011111: finv2 = 23'b11001100000010100010100;
12'b011111100000: finv2 = 23'b11001011111000111010000;
12'b011111100001: finv2 = 23'b11001011101111010001110;
12'b011111100010: finv2 = 23'b11001011100101101001110;
12'b011111100011: finv2 = 23'b11001011011100000010001;
12'b011111100100: finv2 = 23'b11001011010010011010110;
12'b011111100101: finv2 = 23'b11001011001000110011110;
12'b011111100110: finv2 = 23'b11001010111111001101000;
12'b011111100111: finv2 = 23'b11001010110101100110101;
12'b011111101000: finv2 = 23'b11001010101100000000100;
12'b011111101001: finv2 = 23'b11001010100010011010101;
12'b011111101010: finv2 = 23'b11001010011000110101001;
12'b011111101011: finv2 = 23'b11001010001111001111111;
12'b011111101100: finv2 = 23'b11001010000101101010111;
12'b011111101101: finv2 = 23'b11001001111100000110010;
12'b011111101110: finv2 = 23'b11001001110010100010000;
12'b011111101111: finv2 = 23'b11001001101000111101111;
12'b011111110000: finv2 = 23'b11001001011111011010010;
12'b011111110001: finv2 = 23'b11001001010101110110110;
12'b011111110010: finv2 = 23'b11001001001100010011101;
12'b011111110011: finv2 = 23'b11001001000010110000110;
12'b011111110100: finv2 = 23'b11001000111001001110010;
12'b011111110101: finv2 = 23'b11001000101111101100000;
12'b011111110110: finv2 = 23'b11001000100110001010001;
12'b011111110111: finv2 = 23'b11001000011100101000100;
12'b011111111000: finv2 = 23'b11001000010011000111001;
12'b011111111001: finv2 = 23'b11001000001001100110001;
12'b011111111010: finv2 = 23'b11001000000000000101011;
12'b011111111011: finv2 = 23'b11000111110110100100111;
12'b011111111100: finv2 = 23'b11000111101101000100110;
12'b011111111101: finv2 = 23'b11000111100011100100111;
12'b011111111110: finv2 = 23'b11000111011010000101011;
12'b011111111111: finv2 = 23'b11000111010000100110001;
12'b100000000000: finv2 = 23'b11000111000111000111001;
12'b100000000001: finv2 = 23'b11000110111101101000100;
12'b100000000010: finv2 = 23'b11000110110100001010001;
12'b100000000011: finv2 = 23'b11000110101010101100000;
12'b100000000100: finv2 = 23'b11000110100001001110010;
12'b100000000101: finv2 = 23'b11000110010111110000110;
12'b100000000110: finv2 = 23'b11000110001110010011100;
12'b100000000111: finv2 = 23'b11000110000100110110101;
12'b100000001000: finv2 = 23'b11000101111011011010000;
12'b100000001001: finv2 = 23'b11000101110001111101110;
12'b100000001010: finv2 = 23'b11000101101000100001110;
12'b100000001011: finv2 = 23'b11000101011111000110000;
12'b100000001100: finv2 = 23'b11000101010101101010101;
12'b100000001101: finv2 = 23'b11000101001100001111100;
12'b100000001110: finv2 = 23'b11000101000010110100101;
12'b100000001111: finv2 = 23'b11000100111001011010001;
12'b100000010000: finv2 = 23'b11000100101111111111111;
12'b100000010001: finv2 = 23'b11000100100110100101111;
12'b100000010010: finv2 = 23'b11000100011101001100010;
12'b100000010011: finv2 = 23'b11000100010011110010111;
12'b100000010100: finv2 = 23'b11000100001010011001111;
12'b100000010101: finv2 = 23'b11000100000001000001000;
12'b100000010110: finv2 = 23'b11000011110111101000100;
12'b100000010111: finv2 = 23'b11000011101110010000011;
12'b100000011000: finv2 = 23'b11000011100100111000100;
12'b100000011001: finv2 = 23'b11000011011011100000111;
12'b100000011010: finv2 = 23'b11000011010010001001100;
12'b100000011011: finv2 = 23'b11000011001000110010100;
12'b100000011100: finv2 = 23'b11000010111111011011110;
12'b100000011101: finv2 = 23'b11000010110110000101010;
12'b100000011110: finv2 = 23'b11000010101100101111001;
12'b100000011111: finv2 = 23'b11000010100011011001010;
12'b100000100000: finv2 = 23'b11000010011010000011110;
12'b100000100001: finv2 = 23'b11000010010000101110011;
12'b100000100010: finv2 = 23'b11000010000111011001011;
12'b100000100011: finv2 = 23'b11000001111110000100110;
12'b100000100100: finv2 = 23'b11000001110100110000010;
12'b100000100101: finv2 = 23'b11000001101011011100001;
12'b100000100110: finv2 = 23'b11000001100010001000011;
12'b100000100111: finv2 = 23'b11000001011000110100110;
12'b100000101000: finv2 = 23'b11000001001111100001100;
12'b100000101001: finv2 = 23'b11000001000110001110100;
12'b100000101010: finv2 = 23'b11000000111100111011111;
12'b100000101011: finv2 = 23'b11000000110011101001100;
12'b100000101100: finv2 = 23'b11000000101010010111011;
12'b100000101101: finv2 = 23'b11000000100001000101100;
12'b100000101110: finv2 = 23'b11000000010111110100000;
12'b100000101111: finv2 = 23'b11000000001110100010110;
12'b100000110000: finv2 = 23'b11000000000101010001110;
12'b100000110001: finv2 = 23'b10111111111100000001001;
12'b100000110010: finv2 = 23'b10111111110010110000110;
12'b100000110011: finv2 = 23'b10111111101001100000101;
12'b100000110100: finv2 = 23'b10111111100000010000111;
12'b100000110101: finv2 = 23'b10111111010111000001011;
12'b100000110110: finv2 = 23'b10111111001101110010001;
12'b100000110111: finv2 = 23'b10111111000100100011001;
12'b100000111000: finv2 = 23'b10111110111011010100100;
12'b100000111001: finv2 = 23'b10111110110010000110001;
12'b100000111010: finv2 = 23'b10111110101000111000000;
12'b100000111011: finv2 = 23'b10111110011111101010010;
12'b100000111100: finv2 = 23'b10111110010110011100110;
12'b100000111101: finv2 = 23'b10111110001101001111100;
12'b100000111110: finv2 = 23'b10111110000100000010100;
12'b100000111111: finv2 = 23'b10111101111010110101111;
12'b100001000000: finv2 = 23'b10111101110001101001100;
12'b100001000001: finv2 = 23'b10111101101000011101011;
12'b100001000010: finv2 = 23'b10111101011111010001100;
12'b100001000011: finv2 = 23'b10111101010110000110000;
12'b100001000100: finv2 = 23'b10111101001100111010110;
12'b100001000101: finv2 = 23'b10111101000011101111110;
12'b100001000110: finv2 = 23'b10111100111010100101001;
12'b100001000111: finv2 = 23'b10111100110001011010110;
12'b100001001000: finv2 = 23'b10111100101000010000101;
12'b100001001001: finv2 = 23'b10111100011111000110110;
12'b100001001010: finv2 = 23'b10111100010101111101010;
12'b100001001011: finv2 = 23'b10111100001100110100000;
12'b100001001100: finv2 = 23'b10111100000011101011000;
12'b100001001101: finv2 = 23'b10111011111010100010010;
12'b100001001110: finv2 = 23'b10111011110001011001111;
12'b100001001111: finv2 = 23'b10111011101000010001110;
12'b100001010000: finv2 = 23'b10111011011111001001111;
12'b100001010001: finv2 = 23'b10111011010110000010010;
12'b100001010010: finv2 = 23'b10111011001100111011000;
12'b100001010011: finv2 = 23'b10111011000011110100000;
12'b100001010100: finv2 = 23'b10111010111010101101010;
12'b100001010101: finv2 = 23'b10111010110001100110111;
12'b100001010110: finv2 = 23'b10111010101000100000101;
12'b100001010111: finv2 = 23'b10111010011111011010110;
12'b100001011000: finv2 = 23'b10111010010110010101001;
12'b100001011001: finv2 = 23'b10111010001101001111111;
12'b100001011010: finv2 = 23'b10111010000100001010110;
12'b100001011011: finv2 = 23'b10111001111011000110000;
12'b100001011100: finv2 = 23'b10111001110010000001100;
12'b100001011101: finv2 = 23'b10111001101000111101010;
12'b100001011110: finv2 = 23'b10111001011111111001011;
12'b100001011111: finv2 = 23'b10111001010110110101110;
12'b100001100000: finv2 = 23'b10111001001101110010011;
12'b100001100001: finv2 = 23'b10111001000100101111010;
12'b100001100010: finv2 = 23'b10111000111011101100011;
12'b100001100011: finv2 = 23'b10111000110010101001111;
12'b100001100100: finv2 = 23'b10111000101001100111101;
12'b100001100101: finv2 = 23'b10111000100000100101101;
12'b100001100110: finv2 = 23'b10111000010111100011111;
12'b100001100111: finv2 = 23'b10111000001110100010100;
12'b100001101000: finv2 = 23'b10111000000101100001011;
12'b100001101001: finv2 = 23'b10110111111100100000100;
12'b100001101010: finv2 = 23'b10110111110011011111111;
12'b100001101011: finv2 = 23'b10110111101010011111100;
12'b100001101100: finv2 = 23'b10110111100001011111100;
12'b100001101101: finv2 = 23'b10110111011000011111110;
12'b100001101110: finv2 = 23'b10110111001111100000010;
12'b100001101111: finv2 = 23'b10110111000110100001000;
12'b100001110000: finv2 = 23'b10110110111101100010000;
12'b100001110001: finv2 = 23'b10110110110100100011011;
12'b100001110010: finv2 = 23'b10110110101011100101000;
12'b100001110011: finv2 = 23'b10110110100010100110111;
12'b100001110100: finv2 = 23'b10110110011001101001000;
12'b100001110101: finv2 = 23'b10110110010000101011100;
12'b100001110110: finv2 = 23'b10110110000111101110010;
12'b100001110111: finv2 = 23'b10110101111110110001001;
12'b100001111000: finv2 = 23'b10110101110101110100011;
12'b100001111001: finv2 = 23'b10110101101100111000000;
12'b100001111010: finv2 = 23'b10110101100011111011110;
12'b100001111011: finv2 = 23'b10110101011010111111111;
12'b100001111100: finv2 = 23'b10110101010010000100010;
12'b100001111101: finv2 = 23'b10110101001001001000111;
12'b100001111110: finv2 = 23'b10110101000000001101110;
12'b100001111111: finv2 = 23'b10110100110111010010111;
12'b100010000000: finv2 = 23'b10110100101110011000011;
12'b100010000001: finv2 = 23'b10110100100101011110001;
12'b100010000010: finv2 = 23'b10110100011100100100001;
12'b100010000011: finv2 = 23'b10110100010011101010011;
12'b100010000100: finv2 = 23'b10110100001010110000111;
12'b100010000101: finv2 = 23'b10110100000001110111110;
12'b100010000110: finv2 = 23'b10110011111000111110110;
12'b100010000111: finv2 = 23'b10110011110000000110001;
12'b100010001000: finv2 = 23'b10110011100111001101110;
12'b100010001001: finv2 = 23'b10110011011110010101101;
12'b100010001010: finv2 = 23'b10110011010101011101111;
12'b100010001011: finv2 = 23'b10110011001100100110010;
12'b100010001100: finv2 = 23'b10110011000011101111000;
12'b100010001101: finv2 = 23'b10110010111010111000000;
12'b100010001110: finv2 = 23'b10110010110010000001010;
12'b100010001111: finv2 = 23'b10110010101001001010110;
12'b100010010000: finv2 = 23'b10110010100000010100100;
12'b100010010001: finv2 = 23'b10110010010111011110101;
12'b100010010010: finv2 = 23'b10110010001110101000111;
12'b100010010011: finv2 = 23'b10110010000101110011100;
12'b100010010100: finv2 = 23'b10110001111100111110011;
12'b100010010101: finv2 = 23'b10110001110100001001100;
12'b100010010110: finv2 = 23'b10110001101011010100111;
12'b100010010111: finv2 = 23'b10110001100010100000101;
12'b100010011000: finv2 = 23'b10110001011001101100100;
12'b100010011001: finv2 = 23'b10110001010000111000110;
12'b100010011010: finv2 = 23'b10110001001000000101010;
12'b100010011011: finv2 = 23'b10110000111111010010000;
12'b100010011100: finv2 = 23'b10110000110110011111000;
12'b100010011101: finv2 = 23'b10110000101101101100011;
12'b100010011110: finv2 = 23'b10110000100100111001111;
12'b100010011111: finv2 = 23'b10110000011100000111110;
12'b100010100000: finv2 = 23'b10110000010011010101110;
12'b100010100001: finv2 = 23'b10110000001010100100001;
12'b100010100010: finv2 = 23'b10110000000001110010110;
12'b100010100011: finv2 = 23'b10101111111001000001101;
12'b100010100100: finv2 = 23'b10101111110000010000111;
12'b100010100101: finv2 = 23'b10101111100111100000010;
12'b100010100110: finv2 = 23'b10101111011110110000000;
12'b100010100111: finv2 = 23'b10101111010101111111111;
12'b100010101000: finv2 = 23'b10101111001101010000001;
12'b100010101001: finv2 = 23'b10101111000100100000101;
12'b100010101010: finv2 = 23'b10101110111011110001011;
12'b100010101011: finv2 = 23'b10101110110011000010011;
12'b100010101100: finv2 = 23'b10101110101010010011110;
12'b100010101101: finv2 = 23'b10101110100001100101010;
12'b100010101110: finv2 = 23'b10101110011000110111001;
12'b100010101111: finv2 = 23'b10101110010000001001001;
12'b100010110000: finv2 = 23'b10101110000111011011100;
12'b100010110001: finv2 = 23'b10101101111110101110001;
12'b100010110010: finv2 = 23'b10101101110110000001000;
12'b100010110011: finv2 = 23'b10101101101101010100001;
12'b100010110100: finv2 = 23'b10101101100100100111101;
12'b100010110101: finv2 = 23'b10101101011011111011010;
12'b100010110110: finv2 = 23'b10101101010011001111001;
12'b100010110111: finv2 = 23'b10101101001010100011011;
12'b100010111000: finv2 = 23'b10101101000001110111111;
12'b100010111001: finv2 = 23'b10101100111001001100101;
12'b100010111010: finv2 = 23'b10101100110000100001100;
12'b100010111011: finv2 = 23'b10101100100111110110111;
12'b100010111100: finv2 = 23'b10101100011111001100011;
12'b100010111101: finv2 = 23'b10101100010110100010001;
12'b100010111110: finv2 = 23'b10101100001101111000001;
12'b100010111111: finv2 = 23'b10101100000101001110100;
12'b100011000000: finv2 = 23'b10101011111100100101000;
12'b100011000001: finv2 = 23'b10101011110011111011111;
12'b100011000010: finv2 = 23'b10101011101011010010111;
12'b100011000011: finv2 = 23'b10101011100010101010010;
12'b100011000100: finv2 = 23'b10101011011010000001111;
12'b100011000101: finv2 = 23'b10101011010001011001110;
12'b100011000110: finv2 = 23'b10101011001000110001111;
12'b100011000111: finv2 = 23'b10101011000000001010010;
12'b100011001000: finv2 = 23'b10101010110111100011000;
12'b100011001001: finv2 = 23'b10101010101110111011111;
12'b100011001010: finv2 = 23'b10101010100110010101000;
12'b100011001011: finv2 = 23'b10101010011101101110100;
12'b100011001100: finv2 = 23'b10101010010101001000001;
12'b100011001101: finv2 = 23'b10101010001100100010001;
12'b100011001110: finv2 = 23'b10101010000011111100011;
12'b100011001111: finv2 = 23'b10101001111011010110111;
12'b100011010000: finv2 = 23'b10101001110010110001100;
12'b100011010001: finv2 = 23'b10101001101010001100100;
12'b100011010010: finv2 = 23'b10101001100001100111110;
12'b100011010011: finv2 = 23'b10101001011001000011011;
12'b100011010100: finv2 = 23'b10101001010000011111001;
12'b100011010101: finv2 = 23'b10101001000111111011001;
12'b100011010110: finv2 = 23'b10101000111111010111011;
12'b100011010111: finv2 = 23'b10101000110110110100000;
12'b100011011000: finv2 = 23'b10101000101110010000110;
12'b100011011001: finv2 = 23'b10101000100101101101111;
12'b100011011010: finv2 = 23'b10101000011101001011001;
12'b100011011011: finv2 = 23'b10101000010100101000110;
12'b100011011100: finv2 = 23'b10101000001100000110101;
12'b100011011101: finv2 = 23'b10101000000011100100101;
12'b100011011110: finv2 = 23'b10100111111011000011000;
12'b100011011111: finv2 = 23'b10100111110010100001101;
12'b100011100000: finv2 = 23'b10100111101010000000100;
12'b100011100001: finv2 = 23'b10100111100001011111101;
12'b100011100010: finv2 = 23'b10100111011000111111000;
12'b100011100011: finv2 = 23'b10100111010000011110101;
12'b100011100100: finv2 = 23'b10100111000111111110100;
12'b100011100101: finv2 = 23'b10100110111111011110101;
12'b100011100110: finv2 = 23'b10100110110110111111001;
12'b100011100111: finv2 = 23'b10100110101110011111110;
12'b100011101000: finv2 = 23'b10100110100110000000101;
12'b100011101001: finv2 = 23'b10100110011101100001111;
12'b100011101010: finv2 = 23'b10100110010101000011010;
12'b100011101011: finv2 = 23'b10100110001100100101000;
12'b100011101100: finv2 = 23'b10100110000100000110111;
12'b100011101101: finv2 = 23'b10100101111011101001001;
12'b100011101110: finv2 = 23'b10100101110011001011100;
12'b100011101111: finv2 = 23'b10100101101010101110010;
12'b100011110000: finv2 = 23'b10100101100010010001001;
12'b100011110001: finv2 = 23'b10100101011001110100011;
12'b100011110010: finv2 = 23'b10100101010001010111111;
12'b100011110011: finv2 = 23'b10100101001000111011101;
12'b100011110100: finv2 = 23'b10100101000000011111100;
12'b100011110101: finv2 = 23'b10100100111000000011110;
12'b100011110110: finv2 = 23'b10100100101111101000010;
12'b100011110111: finv2 = 23'b10100100100111001101000;
12'b100011111000: finv2 = 23'b10100100011110110010000;
12'b100011111001: finv2 = 23'b10100100010110010111010;
12'b100011111010: finv2 = 23'b10100100001101111100101;
12'b100011111011: finv2 = 23'b10100100000101100010011;
12'b100011111100: finv2 = 23'b10100011111101001000011;
12'b100011111101: finv2 = 23'b10100011110100101110101;
12'b100011111110: finv2 = 23'b10100011101100010101001;
12'b100011111111: finv2 = 23'b10100011100011111011111;
12'b100100000000: finv2 = 23'b10100011011011100010111;
12'b100100000001: finv2 = 23'b10100011010011001010001;
12'b100100000010: finv2 = 23'b10100011001010110001101;
12'b100100000011: finv2 = 23'b10100011000010011001011;
12'b100100000100: finv2 = 23'b10100010111010000001100;
12'b100100000101: finv2 = 23'b10100010110001101001110;
12'b100100000110: finv2 = 23'b10100010101001010010010;
12'b100100000111: finv2 = 23'b10100010100000111011000;
12'b100100001000: finv2 = 23'b10100010011000100100000;
12'b100100001001: finv2 = 23'b10100010010000001101010;
12'b100100001010: finv2 = 23'b10100010000111110110110;
12'b100100001011: finv2 = 23'b10100001111111100000100;
12'b100100001100: finv2 = 23'b10100001110111001010100;
12'b100100001101: finv2 = 23'b10100001101110110100110;
12'b100100001110: finv2 = 23'b10100001100110011111011;
12'b100100001111: finv2 = 23'b10100001011110001010001;
12'b100100010000: finv2 = 23'b10100001010101110101001;
12'b100100010001: finv2 = 23'b10100001001101100000011;
12'b100100010010: finv2 = 23'b10100001000101001011111;
12'b100100010011: finv2 = 23'b10100000111100110111101;
12'b100100010100: finv2 = 23'b10100000110100100011101;
12'b100100010101: finv2 = 23'b10100000101100001111111;
12'b100100010110: finv2 = 23'b10100000100011111100011;
12'b100100010111: finv2 = 23'b10100000011011101001001;
12'b100100011000: finv2 = 23'b10100000010011010110001;
12'b100100011001: finv2 = 23'b10100000001011000011011;
12'b100100011010: finv2 = 23'b10100000000010110000111;
12'b100100011011: finv2 = 23'b10011111111010011110101;
12'b100100011100: finv2 = 23'b10011111110010001100101;
12'b100100011101: finv2 = 23'b10011111101001111010111;
12'b100100011110: finv2 = 23'b10011111100001101001011;
12'b100100011111: finv2 = 23'b10011111011001011000001;
12'b100100100000: finv2 = 23'b10011111010001000111000;
12'b100100100001: finv2 = 23'b10011111001000110110010;
12'b100100100010: finv2 = 23'b10011111000000100101110;
12'b100100100011: finv2 = 23'b10011110111000010101100;
12'b100100100100: finv2 = 23'b10011110110000000101011;
12'b100100100101: finv2 = 23'b10011110100111110101101;
12'b100100100110: finv2 = 23'b10011110011111100110001;
12'b100100100111: finv2 = 23'b10011110010111010110110;
12'b100100101000: finv2 = 23'b10011110001111000111110;
12'b100100101001: finv2 = 23'b10011110000110111000111;
12'b100100101010: finv2 = 23'b10011101111110101010011;
12'b100100101011: finv2 = 23'b10011101110110011100000;
12'b100100101100: finv2 = 23'b10011101101110001110000;
12'b100100101101: finv2 = 23'b10011101100110000000001;
12'b100100101110: finv2 = 23'b10011101011101110010101;
12'b100100101111: finv2 = 23'b10011101010101100101010;
12'b100100110000: finv2 = 23'b10011101001101011000001;
12'b100100110001: finv2 = 23'b10011101000101001011010;
12'b100100110010: finv2 = 23'b10011100111100111110110;
12'b100100110011: finv2 = 23'b10011100110100110010011;
12'b100100110100: finv2 = 23'b10011100101100100110010;
12'b100100110101: finv2 = 23'b10011100100100011010011;
12'b100100110110: finv2 = 23'b10011100011100001110110;
12'b100100110111: finv2 = 23'b10011100010100000011011;
12'b100100111000: finv2 = 23'b10011100001011111000010;
12'b100100111001: finv2 = 23'b10011100000011101101010;
12'b100100111010: finv2 = 23'b10011011111011100010101;
12'b100100111011: finv2 = 23'b10011011110011011000010;
12'b100100111100: finv2 = 23'b10011011101011001110000;
12'b100100111101: finv2 = 23'b10011011100011000100001;
12'b100100111110: finv2 = 23'b10011011011010111010011;
12'b100100111111: finv2 = 23'b10011011010010110001000;
12'b100101000000: finv2 = 23'b10011011001010100111110;
12'b100101000001: finv2 = 23'b10011011000010011110111;
12'b100101000010: finv2 = 23'b10011010111010010110001;
12'b100101000011: finv2 = 23'b10011010110010001101101;
12'b100101000100: finv2 = 23'b10011010101010000101011;
12'b100101000101: finv2 = 23'b10011010100001111101011;
12'b100101000110: finv2 = 23'b10011010011001110101101;
12'b100101000111: finv2 = 23'b10011010010001101110001;
12'b100101001000: finv2 = 23'b10011010001001100110111;
12'b100101001001: finv2 = 23'b10011010000001011111111;
12'b100101001010: finv2 = 23'b10011001111001011001000;
12'b100101001011: finv2 = 23'b10011001110001010010100;
12'b100101001100: finv2 = 23'b10011001101001001100001;
12'b100101001101: finv2 = 23'b10011001100001000110001;
12'b100101001110: finv2 = 23'b10011001011001000000010;
12'b100101001111: finv2 = 23'b10011001010000111010110;
12'b100101010000: finv2 = 23'b10011001001000110101011;
12'b100101010001: finv2 = 23'b10011001000000110000010;
12'b100101010010: finv2 = 23'b10011000111000101011011;
12'b100101010011: finv2 = 23'b10011000110000100110110;
12'b100101010100: finv2 = 23'b10011000101000100010011;
12'b100101010101: finv2 = 23'b10011000100000011110001;
12'b100101010110: finv2 = 23'b10011000011000011010010;
12'b100101010111: finv2 = 23'b10011000010000010110101;
12'b100101011000: finv2 = 23'b10011000001000010011001;
12'b100101011001: finv2 = 23'b10011000000000001111111;
12'b100101011010: finv2 = 23'b10010111111000001101000;
12'b100101011011: finv2 = 23'b10010111110000001010010;
12'b100101011100: finv2 = 23'b10010111101000000111110;
12'b100101011101: finv2 = 23'b10010111100000000101100;
12'b100101011110: finv2 = 23'b10010111011000000011100;
12'b100101011111: finv2 = 23'b10010111010000000001110;
12'b100101100000: finv2 = 23'b10010111001000000000001;
12'b100101100001: finv2 = 23'b10010110111111111110111;
12'b100101100010: finv2 = 23'b10010110110111111101111;
12'b100101100011: finv2 = 23'b10010110101111111101000;
12'b100101100100: finv2 = 23'b10010110100111111100011;
12'b100101100101: finv2 = 23'b10010110011111111100000;
12'b100101100110: finv2 = 23'b10010110010111111011111;
12'b100101100111: finv2 = 23'b10010110001111111100000;
12'b100101101000: finv2 = 23'b10010110000111111100011;
12'b100101101001: finv2 = 23'b10010101111111111101000;
12'b100101101010: finv2 = 23'b10010101110111111101111;
12'b100101101011: finv2 = 23'b10010101101111111110111;
12'b100101101100: finv2 = 23'b10010101101000000000010;
12'b100101101101: finv2 = 23'b10010101100000000001110;
12'b100101101110: finv2 = 23'b10010101011000000011100;
12'b100101101111: finv2 = 23'b10010101010000000101100;
12'b100101110000: finv2 = 23'b10010101001000000111110;
12'b100101110001: finv2 = 23'b10010101000000001010010;
12'b100101110010: finv2 = 23'b10010100111000001100111;
12'b100101110011: finv2 = 23'b10010100110000001111111;
12'b100101110100: finv2 = 23'b10010100101000010011000;
12'b100101110101: finv2 = 23'b10010100100000010110100;
12'b100101110110: finv2 = 23'b10010100011000011010001;
12'b100101110111: finv2 = 23'b10010100010000011110000;
12'b100101111000: finv2 = 23'b10010100001000100010001;
12'b100101111001: finv2 = 23'b10010100000000100110011;
12'b100101111010: finv2 = 23'b10010011111000101011000;
12'b100101111011: finv2 = 23'b10010011110000101111111;
12'b100101111100: finv2 = 23'b10010011101000110100111;
12'b100101111101: finv2 = 23'b10010011100000111010001;
12'b100101111110: finv2 = 23'b10010011011000111111101;
12'b100101111111: finv2 = 23'b10010011010001000101011;
12'b100110000000: finv2 = 23'b10010011001001001011011;
12'b100110000001: finv2 = 23'b10010011000001010001101;
12'b100110000010: finv2 = 23'b10010010111001011000000;
12'b100110000011: finv2 = 23'b10010010110001011110110;
12'b100110000100: finv2 = 23'b10010010101001100101101;
12'b100110000101: finv2 = 23'b10010010100001101100110;
12'b100110000110: finv2 = 23'b10010010011001110100001;
12'b100110000111: finv2 = 23'b10010010010001111011110;
12'b100110001000: finv2 = 23'b10010010001010000011101;
12'b100110001001: finv2 = 23'b10010010000010001011101;
12'b100110001010: finv2 = 23'b10010001111010010100000;
12'b100110001011: finv2 = 23'b10010001110010011100100;
12'b100110001100: finv2 = 23'b10010001101010100101010;
12'b100110001101: finv2 = 23'b10010001100010101110010;
12'b100110001110: finv2 = 23'b10010001011010110111011;
12'b100110001111: finv2 = 23'b10010001010011000000111;
12'b100110010000: finv2 = 23'b10010001001011001010101;
12'b100110010001: finv2 = 23'b10010001000011010100100;
12'b100110010010: finv2 = 23'b10010000111011011110101;
12'b100110010011: finv2 = 23'b10010000110011101001000;
12'b100110010100: finv2 = 23'b10010000101011110011101;
12'b100110010101: finv2 = 23'b10010000100011111110011;
12'b100110010110: finv2 = 23'b10010000011100001001100;
12'b100110010111: finv2 = 23'b10010000010100010100110;
12'b100110011000: finv2 = 23'b10010000001100100000010;
12'b100110011001: finv2 = 23'b10010000000100101100000;
12'b100110011010: finv2 = 23'b10001111111100111000000;
12'b100110011011: finv2 = 23'b10001111110101000100010;
12'b100110011100: finv2 = 23'b10001111101101010000101;
12'b100110011101: finv2 = 23'b10001111100101011101011;
12'b100110011110: finv2 = 23'b10001111011101101010010;
12'b100110011111: finv2 = 23'b10001111010101110111011;
12'b100110100000: finv2 = 23'b10001111001110000100101;
12'b100110100001: finv2 = 23'b10001111000110010010010;
12'b100110100010: finv2 = 23'b10001110111110100000000;
12'b100110100011: finv2 = 23'b10001110110110101110001;
12'b100110100100: finv2 = 23'b10001110101110111100011;
12'b100110100101: finv2 = 23'b10001110100111001010111;
12'b100110100110: finv2 = 23'b10001110011111011001100;
12'b100110100111: finv2 = 23'b10001110010111101000100;
12'b100110101000: finv2 = 23'b10001110001111110111101;
12'b100110101001: finv2 = 23'b10001110001000000111000;
12'b100110101010: finv2 = 23'b10001110000000010110101;
12'b100110101011: finv2 = 23'b10001101111000100110100;
12'b100110101100: finv2 = 23'b10001101110000110110101;
12'b100110101101: finv2 = 23'b10001101101001000110111;
12'b100110101110: finv2 = 23'b10001101100001010111011;
12'b100110101111: finv2 = 23'b10001101011001101000001;
12'b100110110000: finv2 = 23'b10001101010001111001001;
12'b100110110001: finv2 = 23'b10001101001010001010011;
12'b100110110010: finv2 = 23'b10001101000010011011110;
12'b100110110011: finv2 = 23'b10001100111010101101100;
12'b100110110100: finv2 = 23'b10001100110010111111011;
12'b100110110101: finv2 = 23'b10001100101011010001100;
12'b100110110110: finv2 = 23'b10001100100011100011110;
12'b100110110111: finv2 = 23'b10001100011011110110011;
12'b100110111000: finv2 = 23'b10001100010100001001001;
12'b100110111001: finv2 = 23'b10001100001100011100001;
12'b100110111010: finv2 = 23'b10001100000100101111011;
12'b100110111011: finv2 = 23'b10001011111101000010110;
12'b100110111100: finv2 = 23'b10001011110101010110100;
12'b100110111101: finv2 = 23'b10001011101101101010011;
12'b100110111110: finv2 = 23'b10001011100101111110100;
12'b100110111111: finv2 = 23'b10001011011110010010111;
12'b100111000000: finv2 = 23'b10001011010110100111100;
12'b100111000001: finv2 = 23'b10001011001110111100010;
12'b100111000010: finv2 = 23'b10001011000111010001010;
12'b100111000011: finv2 = 23'b10001010111111100110100;
12'b100111000100: finv2 = 23'b10001010110111111100000;
12'b100111000101: finv2 = 23'b10001010110000010001101;
12'b100111000110: finv2 = 23'b10001010101000100111101;
12'b100111000111: finv2 = 23'b10001010100000111101110;
12'b100111001000: finv2 = 23'b10001010011001010100001;
12'b100111001001: finv2 = 23'b10001010010001101010101;
12'b100111001010: finv2 = 23'b10001010001010000001100;
12'b100111001011: finv2 = 23'b10001010000010011000100;
12'b100111001100: finv2 = 23'b10001001111010101111110;
12'b100111001101: finv2 = 23'b10001001110011000111010;
12'b100111001110: finv2 = 23'b10001001101011011110111;
12'b100111001111: finv2 = 23'b10001001100011110110111;
12'b100111010000: finv2 = 23'b10001001011100001111000;
12'b100111010001: finv2 = 23'b10001001010100100111011;
12'b100111010010: finv2 = 23'b10001001001100111111111;
12'b100111010011: finv2 = 23'b10001001000101011000110;
12'b100111010100: finv2 = 23'b10001000111101110001110;
12'b100111010101: finv2 = 23'b10001000110110001011000;
12'b100111010110: finv2 = 23'b10001000101110100100011;
12'b100111010111: finv2 = 23'b10001000100110111110001;
12'b100111011000: finv2 = 23'b10001000011111011000000;
12'b100111011001: finv2 = 23'b10001000010111110010001;
12'b100111011010: finv2 = 23'b10001000010000001100100;
12'b100111011011: finv2 = 23'b10001000001000100111000;
12'b100111011100: finv2 = 23'b10001000000001000001111;
12'b100111011101: finv2 = 23'b10000111111001011100111;
12'b100111011110: finv2 = 23'b10000111110001111000001;
12'b100111011111: finv2 = 23'b10000111101010010011100;
12'b100111100000: finv2 = 23'b10000111100010101111001;
12'b100111100001: finv2 = 23'b10000111011011001011000;
12'b100111100010: finv2 = 23'b10000111010011100111001;
12'b100111100011: finv2 = 23'b10000111001100000011100;
12'b100111100100: finv2 = 23'b10000111000100100000000;
12'b100111100101: finv2 = 23'b10000110111100111100110;
12'b100111100110: finv2 = 23'b10000110110101011001110;
12'b100111100111: finv2 = 23'b10000110101101110111000;
12'b100111101000: finv2 = 23'b10000110100110010100011;
12'b100111101001: finv2 = 23'b10000110011110110010000;
12'b100111101010: finv2 = 23'b10000110010111001111111;
12'b100111101011: finv2 = 23'b10000110001111101101111;
12'b100111101100: finv2 = 23'b10000110001000001100010;
12'b100111101101: finv2 = 23'b10000110000000101010110;
12'b100111101110: finv2 = 23'b10000101111001001001011;
12'b100111101111: finv2 = 23'b10000101110001101000011;
12'b100111110000: finv2 = 23'b10000101101010000111100;
12'b100111110001: finv2 = 23'b10000101100010100110111;
12'b100111110010: finv2 = 23'b10000101011011000110100;
12'b100111110011: finv2 = 23'b10000101010011100110010;
12'b100111110100: finv2 = 23'b10000101001100000110011;
12'b100111110101: finv2 = 23'b10000101000100100110100;
12'b100111110110: finv2 = 23'b10000100111101000111000;
12'b100111110111: finv2 = 23'b10000100110101100111110;
12'b100111111000: finv2 = 23'b10000100101110001000101;
12'b100111111001: finv2 = 23'b10000100100110101001110;
12'b100111111010: finv2 = 23'b10000100011111001011000;
12'b100111111011: finv2 = 23'b10000100010111101100100;
12'b100111111100: finv2 = 23'b10000100010000001110010;
12'b100111111101: finv2 = 23'b10000100001000110000010;
12'b100111111110: finv2 = 23'b10000100000001010010100;
12'b100111111111: finv2 = 23'b10000011111001110100111;
12'b101000000000: finv2 = 23'b10000011110010010111100;
12'b101000000001: finv2 = 23'b10000011101010111010010;
12'b101000000010: finv2 = 23'b10000011100011011101011;
12'b101000000011: finv2 = 23'b10000011011100000000101;
12'b101000000100: finv2 = 23'b10000011010100100100001;
12'b101000000101: finv2 = 23'b10000011001101000111110;
12'b101000000110: finv2 = 23'b10000011000101101011110;
12'b101000000111: finv2 = 23'b10000010111110001111110;
12'b101000001000: finv2 = 23'b10000010110110110100001;
12'b101000001001: finv2 = 23'b10000010101111011000110;
12'b101000001010: finv2 = 23'b10000010100111111101100;
12'b101000001011: finv2 = 23'b10000010100000100010011;
12'b101000001100: finv2 = 23'b10000010011001000111101;
12'b101000001101: finv2 = 23'b10000010010001101101000;
12'b101000001110: finv2 = 23'b10000010001010010010101;
12'b101000001111: finv2 = 23'b10000010000010111000100;
12'b101000010000: finv2 = 23'b10000001111011011110100;
12'b101000010001: finv2 = 23'b10000001110100000100110;
12'b101000010010: finv2 = 23'b10000001101100101011010;
12'b101000010011: finv2 = 23'b10000001100101010001111;
12'b101000010100: finv2 = 23'b10000001011101111000110;
12'b101000010101: finv2 = 23'b10000001010110011111111;
12'b101000010110: finv2 = 23'b10000001001111000111010;
12'b101000010111: finv2 = 23'b10000001000111101110110;
12'b101000011000: finv2 = 23'b10000001000000010110100;
12'b101000011001: finv2 = 23'b10000000111000111110100;
12'b101000011010: finv2 = 23'b10000000110001100110101;
12'b101000011011: finv2 = 23'b10000000101010001111000;
12'b101000011100: finv2 = 23'b10000000100010110111101;
12'b101000011101: finv2 = 23'b10000000011011100000011;
12'b101000011110: finv2 = 23'b10000000010100001001011;
12'b101000011111: finv2 = 23'b10000000001100110010101;
12'b101000100000: finv2 = 23'b10000000000101011100001;
12'b101000100001: finv2 = 23'b01111111111110000101110;
12'b101000100010: finv2 = 23'b01111111110110101111101;
12'b101000100011: finv2 = 23'b01111111101111011001101;
12'b101000100100: finv2 = 23'b01111111101000000011111;
12'b101000100101: finv2 = 23'b01111111100000101110011;
12'b101000100110: finv2 = 23'b01111111011001011001001;
12'b101000100111: finv2 = 23'b01111111010010000100000;
12'b101000101000: finv2 = 23'b01111111001010101111001;
12'b101000101001: finv2 = 23'b01111111000011011010100;
12'b101000101010: finv2 = 23'b01111110111100000110000;
12'b101000101011: finv2 = 23'b01111110110100110001110;
12'b101000101100: finv2 = 23'b01111110101101011101110;
12'b101000101101: finv2 = 23'b01111110100110001001111;
12'b101000101110: finv2 = 23'b01111110011110110110010;
12'b101000101111: finv2 = 23'b01111110010111100010111;
12'b101000110000: finv2 = 23'b01111110010000001111101;
12'b101000110001: finv2 = 23'b01111110001000111100101;
12'b101000110010: finv2 = 23'b01111110000001101001111;
12'b101000110011: finv2 = 23'b01111101111010010111011;
12'b101000110100: finv2 = 23'b01111101110011000101000;
12'b101000110101: finv2 = 23'b01111101101011110010110;
12'b101000110110: finv2 = 23'b01111101100100100000111;
12'b101000110111: finv2 = 23'b01111101011101001111001;
12'b101000111000: finv2 = 23'b01111101010101111101101;
12'b101000111001: finv2 = 23'b01111101001110101100010;
12'b101000111010: finv2 = 23'b01111101000111011011001;
12'b101000111011: finv2 = 23'b01111101000000001010010;
12'b101000111100: finv2 = 23'b01111100111000111001100;
12'b101000111101: finv2 = 23'b01111100110001101001000;
12'b101000111110: finv2 = 23'b01111100101010011000110;
12'b101000111111: finv2 = 23'b01111100100011001000101;
12'b101001000000: finv2 = 23'b01111100011011111000110;
12'b101001000001: finv2 = 23'b01111100010100101001001;
12'b101001000010: finv2 = 23'b01111100001101011001101;
12'b101001000011: finv2 = 23'b01111100000110001010011;
12'b101001000100: finv2 = 23'b01111011111110111011011;
12'b101001000101: finv2 = 23'b01111011110111101100100;
12'b101001000110: finv2 = 23'b01111011110000011101111;
12'b101001000111: finv2 = 23'b01111011101001001111100;
12'b101001001000: finv2 = 23'b01111011100010000001010;
12'b101001001001: finv2 = 23'b01111011011010110011010;
12'b101001001010: finv2 = 23'b01111011010011100101011;
12'b101001001011: finv2 = 23'b01111011001100010111111;
12'b101001001100: finv2 = 23'b01111011000101001010011;
12'b101001001101: finv2 = 23'b01111010111101111101010;
12'b101001001110: finv2 = 23'b01111010110110110000010;
12'b101001001111: finv2 = 23'b01111010101111100011100;
12'b101001010000: finv2 = 23'b01111010101000010110111;
12'b101001010001: finv2 = 23'b01111010100001001010100;
12'b101001010010: finv2 = 23'b01111010011001111110011;
12'b101001010011: finv2 = 23'b01111010010010110010011;
12'b101001010100: finv2 = 23'b01111010001011100110101;
12'b101001010101: finv2 = 23'b01111010000100011011001;
12'b101001010110: finv2 = 23'b01111001111101001111110;
12'b101001010111: finv2 = 23'b01111001110110000100101;
12'b101001011000: finv2 = 23'b01111001101110111001101;
12'b101001011001: finv2 = 23'b01111001100111101110111;
12'b101001011010: finv2 = 23'b01111001100000100100011;
12'b101001011011: finv2 = 23'b01111001011001011010001;
12'b101001011100: finv2 = 23'b01111001010010010000000;
12'b101001011101: finv2 = 23'b01111001001011000110000;
12'b101001011110: finv2 = 23'b01111001000011111100011;
12'b101001011111: finv2 = 23'b01111000111100110010110;
12'b101001100000: finv2 = 23'b01111000110101101001100;
12'b101001100001: finv2 = 23'b01111000101110100000011;
12'b101001100010: finv2 = 23'b01111000100111010111100;
12'b101001100011: finv2 = 23'b01111000100000001110110;
12'b101001100100: finv2 = 23'b01111000011001000110010;
12'b101001100101: finv2 = 23'b01111000010001111110000;
12'b101001100110: finv2 = 23'b01111000001010110101111;
12'b101001100111: finv2 = 23'b01111000000011101110000;
12'b101001101000: finv2 = 23'b01110111111100100110011;
12'b101001101001: finv2 = 23'b01110111110101011110111;
12'b101001101010: finv2 = 23'b01110111101110010111101;
12'b101001101011: finv2 = 23'b01110111100111010000100;
12'b101001101100: finv2 = 23'b01110111100000001001101;
12'b101001101101: finv2 = 23'b01110111011001000010111;
12'b101001101110: finv2 = 23'b01110111010001111100100;
12'b101001101111: finv2 = 23'b01110111001010110110001;
12'b101001110000: finv2 = 23'b01110111000011110000001;
12'b101001110001: finv2 = 23'b01110110111100101010010;
12'b101001110010: finv2 = 23'b01110110110101100100101;
12'b101001110011: finv2 = 23'b01110110101110011111001;
12'b101001110100: finv2 = 23'b01110110100111011001111;
12'b101001110101: finv2 = 23'b01110110100000010100110;
12'b101001110110: finv2 = 23'b01110110011001001111111;
12'b101001110111: finv2 = 23'b01110110010010001011010;
12'b101001111000: finv2 = 23'b01110110001011000110110;
12'b101001111001: finv2 = 23'b01110110000100000010100;
12'b101001111010: finv2 = 23'b01110101111100111110011;
12'b101001111011: finv2 = 23'b01110101110101111010101;
12'b101001111100: finv2 = 23'b01110101101110110110111;
12'b101001111101: finv2 = 23'b01110101100111110011100;
12'b101001111110: finv2 = 23'b01110101100000110000001;
12'b101001111111: finv2 = 23'b01110101011001101101001;
12'b101010000000: finv2 = 23'b01110101010010101010010;
12'b101010000001: finv2 = 23'b01110101001011100111101;
12'b101010000010: finv2 = 23'b01110101000100100101001;
12'b101010000011: finv2 = 23'b01110100111101100010111;
12'b101010000100: finv2 = 23'b01110100110110100000110;
12'b101010000101: finv2 = 23'b01110100101111011110111;
12'b101010000110: finv2 = 23'b01110100101000011101010;
12'b101010000111: finv2 = 23'b01110100100001011011110;
12'b101010001000: finv2 = 23'b01110100011010011010100;
12'b101010001001: finv2 = 23'b01110100010011011001011;
12'b101010001010: finv2 = 23'b01110100001100011000100;
12'b101010001011: finv2 = 23'b01110100000101010111111;
12'b101010001100: finv2 = 23'b01110011111110010111011;
12'b101010001101: finv2 = 23'b01110011110111010111001;
12'b101010001110: finv2 = 23'b01110011110000010111000;
12'b101010001111: finv2 = 23'b01110011101001010111001;
12'b101010010000: finv2 = 23'b01110011100010010111011;
12'b101010010001: finv2 = 23'b01110011011011010111111;
12'b101010010010: finv2 = 23'b01110011010100011000101;
12'b101010010011: finv2 = 23'b01110011001101011001100;
12'b101010010100: finv2 = 23'b01110011000110011010101;
12'b101010010101: finv2 = 23'b01110010111111011011111;
12'b101010010110: finv2 = 23'b01110010111000011101011;
12'b101010010111: finv2 = 23'b01110010110001011111001;
12'b101010011000: finv2 = 23'b01110010101010100001000;
12'b101010011001: finv2 = 23'b01110010100011100011000;
12'b101010011010: finv2 = 23'b01110010011100100101011;
12'b101010011011: finv2 = 23'b01110010010101100111110;
12'b101010011100: finv2 = 23'b01110010001110101010100;
12'b101010011101: finv2 = 23'b01110010000111101101011;
12'b101010011110: finv2 = 23'b01110010000000110000011;
12'b101010011111: finv2 = 23'b01110001111001110011101;
12'b101010100000: finv2 = 23'b01110001110010110111001;
12'b101010100001: finv2 = 23'b01110001101011111010110;
12'b101010100010: finv2 = 23'b01110001100100111110101;
12'b101010100011: finv2 = 23'b01110001011110000010101;
12'b101010100100: finv2 = 23'b01110001010111000110111;
12'b101010100101: finv2 = 23'b01110001010000001011011;
12'b101010100110: finv2 = 23'b01110001001001010000000;
12'b101010100111: finv2 = 23'b01110001000010010100110;
12'b101010101000: finv2 = 23'b01110000111011011001110;
12'b101010101001: finv2 = 23'b01110000110100011111000;
12'b101010101010: finv2 = 23'b01110000101101100100011;
12'b101010101011: finv2 = 23'b01110000100110101010000;
12'b101010101100: finv2 = 23'b01110000011111101111110;
12'b101010101101: finv2 = 23'b01110000011000110101110;
12'b101010101110: finv2 = 23'b01110000010001111100000;
12'b101010101111: finv2 = 23'b01110000001011000010011;
12'b101010110000: finv2 = 23'b01110000000100001000111;
12'b101010110001: finv2 = 23'b01101111111101001111101;
12'b101010110010: finv2 = 23'b01101111110110010110101;
12'b101010110011: finv2 = 23'b01101111101111011101110;
12'b101010110100: finv2 = 23'b01101111101000100101001;
12'b101010110101: finv2 = 23'b01101111100001101100101;
12'b101010110110: finv2 = 23'b01101111011010110100011;
12'b101010110111: finv2 = 23'b01101111010011111100011;
12'b101010111000: finv2 = 23'b01101111001101000100011;
12'b101010111001: finv2 = 23'b01101111000110001100110;
12'b101010111010: finv2 = 23'b01101110111111010101010;
12'b101010111011: finv2 = 23'b01101110111000011110000;
12'b101010111100: finv2 = 23'b01101110110001100110111;
12'b101010111101: finv2 = 23'b01101110101010101111111;
12'b101010111110: finv2 = 23'b01101110100011111001001;
12'b101010111111: finv2 = 23'b01101110011101000010101;
12'b101011000000: finv2 = 23'b01101110010110001100010;
12'b101011000001: finv2 = 23'b01101110001111010110001;
12'b101011000010: finv2 = 23'b01101110001000100000010;
12'b101011000011: finv2 = 23'b01101110000001101010011;
12'b101011000100: finv2 = 23'b01101101111010110100111;
12'b101011000101: finv2 = 23'b01101101110011111111100;
12'b101011000110: finv2 = 23'b01101101101101001010010;
12'b101011000111: finv2 = 23'b01101101100110010101010;
12'b101011001000: finv2 = 23'b01101101011111100000100;
12'b101011001001: finv2 = 23'b01101101011000101011111;
12'b101011001010: finv2 = 23'b01101101010001110111011;
12'b101011001011: finv2 = 23'b01101101001011000011001;
12'b101011001100: finv2 = 23'b01101101000100001111001;
12'b101011001101: finv2 = 23'b01101100111101011011010;
12'b101011001110: finv2 = 23'b01101100110110100111101;
12'b101011001111: finv2 = 23'b01101100101111110100001;
12'b101011010000: finv2 = 23'b01101100101001000000111;
12'b101011010001: finv2 = 23'b01101100100010001101110;
12'b101011010010: finv2 = 23'b01101100011011011010111;
12'b101011010011: finv2 = 23'b01101100010100101000001;
12'b101011010100: finv2 = 23'b01101100001101110101101;
12'b101011010101: finv2 = 23'b01101100000111000011010;
12'b101011010110: finv2 = 23'b01101100000000010001001;
12'b101011010111: finv2 = 23'b01101011111001011111010;
12'b101011011000: finv2 = 23'b01101011110010101101011;
12'b101011011001: finv2 = 23'b01101011101011111011111;
12'b101011011010: finv2 = 23'b01101011100101001010100;
12'b101011011011: finv2 = 23'b01101011011110011001010;
12'b101011011100: finv2 = 23'b01101011010111101000010;
12'b101011011101: finv2 = 23'b01101011010000110111011;
12'b101011011110: finv2 = 23'b01101011001010000110110;
12'b101011011111: finv2 = 23'b01101011000011010110011;
12'b101011100000: finv2 = 23'b01101010111100100110001;
12'b101011100001: finv2 = 23'b01101010110101110110000;
12'b101011100010: finv2 = 23'b01101010101111000110001;
12'b101011100011: finv2 = 23'b01101010101000010110100;
12'b101011100100: finv2 = 23'b01101010100001100111000;
12'b101011100101: finv2 = 23'b01101010011010110111101;
12'b101011100110: finv2 = 23'b01101010010100001000100;
12'b101011100111: finv2 = 23'b01101010001101011001101;
12'b101011101000: finv2 = 23'b01101010000110101010111;
12'b101011101001: finv2 = 23'b01101001111111111100010;
12'b101011101010: finv2 = 23'b01101001111001001101111;
12'b101011101011: finv2 = 23'b01101001110010011111110;
12'b101011101100: finv2 = 23'b01101001101011110001110;
12'b101011101101: finv2 = 23'b01101001100101000011111;
12'b101011101110: finv2 = 23'b01101001011110010110010;
12'b101011101111: finv2 = 23'b01101001010111101000111;
12'b101011110000: finv2 = 23'b01101001010000111011101;
12'b101011110001: finv2 = 23'b01101001001010001110100;
12'b101011110010: finv2 = 23'b01101001000011100001101;
12'b101011110011: finv2 = 23'b01101000111100110101000;
12'b101011110100: finv2 = 23'b01101000110110001000100;
12'b101011110101: finv2 = 23'b01101000101111011100001;
12'b101011110110: finv2 = 23'b01101000101000110000000;
12'b101011110111: finv2 = 23'b01101000100010000100000;
12'b101011111000: finv2 = 23'b01101000011011011000010;
12'b101011111001: finv2 = 23'b01101000010100101100110;
12'b101011111010: finv2 = 23'b01101000001110000001011;
12'b101011111011: finv2 = 23'b01101000000111010110001;
12'b101011111100: finv2 = 23'b01101000000000101011001;
12'b101011111101: finv2 = 23'b01100111111010000000010;
12'b101011111110: finv2 = 23'b01100111110011010101101;
12'b101011111111: finv2 = 23'b01100111101100101011001;
12'b101100000000: finv2 = 23'b01100111100110000000111;
12'b101100000001: finv2 = 23'b01100111011111010110110;
12'b101100000010: finv2 = 23'b01100111011000101100111;
12'b101100000011: finv2 = 23'b01100111010010000011001;
12'b101100000100: finv2 = 23'b01100111001011011001101;
12'b101100000101: finv2 = 23'b01100111000100110000010;
12'b101100000110: finv2 = 23'b01100110111110000111001;
12'b101100000111: finv2 = 23'b01100110110111011110001;
12'b101100001000: finv2 = 23'b01100110110000110101010;
12'b101100001001: finv2 = 23'b01100110101010001100110;
12'b101100001010: finv2 = 23'b01100110100011100100010;
12'b101100001011: finv2 = 23'b01100110011100111100000;
12'b101100001100: finv2 = 23'b01100110010110010100000;
12'b101100001101: finv2 = 23'b01100110001111101100000;
12'b101100001110: finv2 = 23'b01100110001001000100011;
12'b101100001111: finv2 = 23'b01100110000010011100111;
12'b101100010000: finv2 = 23'b01100101111011110101100;
12'b101100010001: finv2 = 23'b01100101110101001110011;
12'b101100010010: finv2 = 23'b01100101101110100111011;
12'b101100010011: finv2 = 23'b01100101101000000000101;
12'b101100010100: finv2 = 23'b01100101100001011010000;
12'b101100010101: finv2 = 23'b01100101011010110011101;
12'b101100010110: finv2 = 23'b01100101010100001101011;
12'b101100010111: finv2 = 23'b01100101001101100111011;
12'b101100011000: finv2 = 23'b01100101000111000001100;
12'b101100011001: finv2 = 23'b01100101000000011011110;
12'b101100011010: finv2 = 23'b01100100111001110110010;
12'b101100011011: finv2 = 23'b01100100110011010001000;
12'b101100011100: finv2 = 23'b01100100101100101011110;
12'b101100011101: finv2 = 23'b01100100100110000110111;
12'b101100011110: finv2 = 23'b01100100011111100010001;
12'b101100011111: finv2 = 23'b01100100011000111101100;
12'b101100100000: finv2 = 23'b01100100010010011001001;
12'b101100100001: finv2 = 23'b01100100001011110100111;
12'b101100100010: finv2 = 23'b01100100000101010000110;
12'b101100100011: finv2 = 23'b01100011111110101100111;
12'b101100100100: finv2 = 23'b01100011111000001001010;
12'b101100100101: finv2 = 23'b01100011110001100101110;
12'b101100100110: finv2 = 23'b01100011101011000010011;
12'b101100100111: finv2 = 23'b01100011100100011111010;
12'b101100101000: finv2 = 23'b01100011011101111100010;
12'b101100101001: finv2 = 23'b01100011010111011001100;
12'b101100101010: finv2 = 23'b01100011010000110110111;
12'b101100101011: finv2 = 23'b01100011001010010100100;
12'b101100101100: finv2 = 23'b01100011000011110010010;
12'b101100101101: finv2 = 23'b01100010111101010000010;
12'b101100101110: finv2 = 23'b01100010110110101110011;
12'b101100101111: finv2 = 23'b01100010110000001100101;
12'b101100110000: finv2 = 23'b01100010101001101011001;
12'b101100110001: finv2 = 23'b01100010100011001001110;
12'b101100110010: finv2 = 23'b01100010011100101000101;
12'b101100110011: finv2 = 23'b01100010010110000111101;
12'b101100110100: finv2 = 23'b01100010001111100110111;
12'b101100110101: finv2 = 23'b01100010001001000110010;
12'b101100110110: finv2 = 23'b01100010000010100101110;
12'b101100110111: finv2 = 23'b01100001111100000101100;
12'b101100111000: finv2 = 23'b01100001110101100101011;
12'b101100111001: finv2 = 23'b01100001101111000101100;
12'b101100111010: finv2 = 23'b01100001101000100101110;
12'b101100111011: finv2 = 23'b01100001100010000110010;
12'b101100111100: finv2 = 23'b01100001011011100110111;
12'b101100111101: finv2 = 23'b01100001010101000111110;
12'b101100111110: finv2 = 23'b01100001001110101000110;
12'b101100111111: finv2 = 23'b01100001001000001001111;
12'b101101000000: finv2 = 23'b01100001000001101011010;
12'b101101000001: finv2 = 23'b01100000111011001100110;
12'b101101000010: finv2 = 23'b01100000110100101110100;
12'b101101000011: finv2 = 23'b01100000101110010000011;
12'b101101000100: finv2 = 23'b01100000100111110010011;
12'b101101000101: finv2 = 23'b01100000100001010100101;
12'b101101000110: finv2 = 23'b01100000011010110111000;
12'b101101000111: finv2 = 23'b01100000010100011001101;
12'b101101001000: finv2 = 23'b01100000001101111100011;
12'b101101001001: finv2 = 23'b01100000000111011111011;
12'b101101001010: finv2 = 23'b01100000000001000010100;
12'b101101001011: finv2 = 23'b01011111111010100101110;
12'b101101001100: finv2 = 23'b01011111110100001001010;
12'b101101001101: finv2 = 23'b01011111101101101100111;
12'b101101001110: finv2 = 23'b01011111100111010000110;
12'b101101001111: finv2 = 23'b01011111100000110100110;
12'b101101010000: finv2 = 23'b01011111011010011001000;
12'b101101010001: finv2 = 23'b01011111010011111101011;
12'b101101010010: finv2 = 23'b01011111001101100001111;
12'b101101010011: finv2 = 23'b01011111000111000110101;
12'b101101010100: finv2 = 23'b01011111000000101011100;
12'b101101010101: finv2 = 23'b01011110111010010000100;
12'b101101010110: finv2 = 23'b01011110110011110101110;
12'b101101010111: finv2 = 23'b01011110101101011011010;
12'b101101011000: finv2 = 23'b01011110100111000000111;
12'b101101011001: finv2 = 23'b01011110100000100110101;
12'b101101011010: finv2 = 23'b01011110011010001100100;
12'b101101011011: finv2 = 23'b01011110010011110010101;
12'b101101011100: finv2 = 23'b01011110001101011001000;
12'b101101011101: finv2 = 23'b01011110000110111111100;
12'b101101011110: finv2 = 23'b01011110000000100110001;
12'b101101011111: finv2 = 23'b01011101111010001100111;
12'b101101100000: finv2 = 23'b01011101110011110011111;
12'b101101100001: finv2 = 23'b01011101101101011011001;
12'b101101100010: finv2 = 23'b01011101100111000010100;
12'b101101100011: finv2 = 23'b01011101100000101010000;
12'b101101100100: finv2 = 23'b01011101011010010001110;
12'b101101100101: finv2 = 23'b01011101010011111001101;
12'b101101100110: finv2 = 23'b01011101001101100001101;
12'b101101100111: finv2 = 23'b01011101000111001001111;
12'b101101101000: finv2 = 23'b01011101000000110010010;
12'b101101101001: finv2 = 23'b01011100111010011010111;
12'b101101101010: finv2 = 23'b01011100110100000011101;
12'b101101101011: finv2 = 23'b01011100101101101100100;
12'b101101101100: finv2 = 23'b01011100100111010101101;
12'b101101101101: finv2 = 23'b01011100100000111110111;
12'b101101101110: finv2 = 23'b01011100011010101000010;
12'b101101101111: finv2 = 23'b01011100010100010001111;
12'b101101110000: finv2 = 23'b01011100001101111011110;
12'b101101110001: finv2 = 23'b01011100000111100101101;
12'b101101110010: finv2 = 23'b01011100000001001111111;
12'b101101110011: finv2 = 23'b01011011111010111010001;
12'b101101110100: finv2 = 23'b01011011110100100100101;
12'b101101110101: finv2 = 23'b01011011101110001111010;
12'b101101110110: finv2 = 23'b01011011100111111010001;
12'b101101110111: finv2 = 23'b01011011100001100101001;
12'b101101111000: finv2 = 23'b01011011011011010000010;
12'b101101111001: finv2 = 23'b01011011010100111011101;
12'b101101111010: finv2 = 23'b01011011001110100111001;
12'b101101111011: finv2 = 23'b01011011001000010010111;
12'b101101111100: finv2 = 23'b01011011000001111110110;
12'b101101111101: finv2 = 23'b01011010111011101010110;
12'b101101111110: finv2 = 23'b01011010110101010111000;
12'b101101111111: finv2 = 23'b01011010101111000011011;
12'b101110000000: finv2 = 23'b01011010101000101111111;
12'b101110000001: finv2 = 23'b01011010100010011100101;
12'b101110000010: finv2 = 23'b01011010011100001001100;
12'b101110000011: finv2 = 23'b01011010010101110110101;
12'b101110000100: finv2 = 23'b01011010001111100011111;
12'b101110000101: finv2 = 23'b01011010001001010001010;
12'b101110000110: finv2 = 23'b01011010000010111110111;
12'b101110000111: finv2 = 23'b01011001111100101100101;
12'b101110001000: finv2 = 23'b01011001110110011010100;
12'b101110001001: finv2 = 23'b01011001110000001000101;
12'b101110001010: finv2 = 23'b01011001101001110110111;
12'b101110001011: finv2 = 23'b01011001100011100101011;
12'b101110001100: finv2 = 23'b01011001011101010100000;
12'b101110001101: finv2 = 23'b01011001010111000010110;
12'b101110001110: finv2 = 23'b01011001010000110001101;
12'b101110001111: finv2 = 23'b01011001001010100000110;
12'b101110010000: finv2 = 23'b01011001000100010000001;
12'b101110010001: finv2 = 23'b01011000111101111111100;
12'b101110010010: finv2 = 23'b01011000110111101111001;
12'b101110010011: finv2 = 23'b01011000110001011111000;
12'b101110010100: finv2 = 23'b01011000101011001111000;
12'b101110010101: finv2 = 23'b01011000100100111111001;
12'b101110010110: finv2 = 23'b01011000011110101111011;
12'b101110010111: finv2 = 23'b01011000011000011111111;
12'b101110011000: finv2 = 23'b01011000010010010000100;
12'b101110011001: finv2 = 23'b01011000001100000001011;
12'b101110011010: finv2 = 23'b01011000000101110010011;
12'b101110011011: finv2 = 23'b01010111111111100011100;
12'b101110011100: finv2 = 23'b01010111111001010100111;
12'b101110011101: finv2 = 23'b01010111110011000110011;
12'b101110011110: finv2 = 23'b01010111101100111000000;
12'b101110011111: finv2 = 23'b01010111100110101001111;
12'b101110100000: finv2 = 23'b01010111100000011011111;
12'b101110100001: finv2 = 23'b01010111011010001110000;
12'b101110100010: finv2 = 23'b01010111010100000000011;
12'b101110100011: finv2 = 23'b01010111001101110010111;
12'b101110100100: finv2 = 23'b01010111000111100101101;
12'b101110100101: finv2 = 23'b01010111000001011000100;
12'b101110100110: finv2 = 23'b01010110111011001011100;
12'b101110100111: finv2 = 23'b01010110110100111110101;
12'b101110101000: finv2 = 23'b01010110101110110010000;
12'b101110101001: finv2 = 23'b01010110101000100101100;
12'b101110101010: finv2 = 23'b01010110100010011001010;
12'b101110101011: finv2 = 23'b01010110011100001101001;
12'b101110101100: finv2 = 23'b01010110010110000001001;
12'b101110101101: finv2 = 23'b01010110001111110101010;
12'b101110101110: finv2 = 23'b01010110001001101001101;
12'b101110101111: finv2 = 23'b01010110000011011110010;
12'b101110110000: finv2 = 23'b01010101111101010010111;
12'b101110110001: finv2 = 23'b01010101110111000111110;
12'b101110110010: finv2 = 23'b01010101110000111100110;
12'b101110110011: finv2 = 23'b01010101101010110010000;
12'b101110110100: finv2 = 23'b01010101100100100111011;
12'b101110110101: finv2 = 23'b01010101011110011100111;
12'b101110110110: finv2 = 23'b01010101011000010010101;
12'b101110110111: finv2 = 23'b01010101010010001000100;
12'b101110111000: finv2 = 23'b01010101001011111110100;
12'b101110111001: finv2 = 23'b01010101000101110100101;
12'b101110111010: finv2 = 23'b01010100111111101011000;
12'b101110111011: finv2 = 23'b01010100111001100001101;
12'b101110111100: finv2 = 23'b01010100110011011000010;
12'b101110111101: finv2 = 23'b01010100101101001111001;
12'b101110111110: finv2 = 23'b01010100100111000110001;
12'b101110111111: finv2 = 23'b01010100100000111101011;
12'b101111000000: finv2 = 23'b01010100011010110100110;
12'b101111000001: finv2 = 23'b01010100010100101100010;
12'b101111000010: finv2 = 23'b01010100001110100100000;
12'b101111000011: finv2 = 23'b01010100001000011011110;
12'b101111000100: finv2 = 23'b01010100000010010011111;
12'b101111000101: finv2 = 23'b01010011111100001100000;
12'b101111000110: finv2 = 23'b01010011110110000100011;
12'b101111000111: finv2 = 23'b01010011101111111100111;
12'b101111001000: finv2 = 23'b01010011101001110101101;
12'b101111001001: finv2 = 23'b01010011100011101110011;
12'b101111001010: finv2 = 23'b01010011011101100111100;
12'b101111001011: finv2 = 23'b01010011010111100000101;
12'b101111001100: finv2 = 23'b01010011010001011010000;
12'b101111001101: finv2 = 23'b01010011001011010011100;
12'b101111001110: finv2 = 23'b01010011000101001101001;
12'b101111001111: finv2 = 23'b01010010111111000111000;
12'b101111010000: finv2 = 23'b01010010111001000001000;
12'b101111010001: finv2 = 23'b01010010110010111011001;
12'b101111010010: finv2 = 23'b01010010101100110101100;
12'b101111010011: finv2 = 23'b01010010100110110000000;
12'b101111010100: finv2 = 23'b01010010100000101010101;
12'b101111010101: finv2 = 23'b01010010011010100101100;
12'b101111010110: finv2 = 23'b01010010010100100000100;
12'b101111010111: finv2 = 23'b01010010001110011011101;
12'b101111011000: finv2 = 23'b01010010001000010110111;
12'b101111011001: finv2 = 23'b01010010000010010010011;
12'b101111011010: finv2 = 23'b01010001111100001110000;
12'b101111011011: finv2 = 23'b01010001110110001001111;
12'b101111011100: finv2 = 23'b01010001110000000101111;
12'b101111011101: finv2 = 23'b01010001101010000010000;
12'b101111011110: finv2 = 23'b01010001100011111110010;
12'b101111011111: finv2 = 23'b01010001011101111010110;
12'b101111100000: finv2 = 23'b01010001010111110111011;
12'b101111100001: finv2 = 23'b01010001010001110100001;
12'b101111100010: finv2 = 23'b01010001001011110001000;
12'b101111100011: finv2 = 23'b01010001000101101110001;
12'b101111100100: finv2 = 23'b01010000111111101011011;
12'b101111100101: finv2 = 23'b01010000111001101000111;
12'b101111100110: finv2 = 23'b01010000110011100110100;
12'b101111100111: finv2 = 23'b01010000101101100100010;
12'b101111101000: finv2 = 23'b01010000100111100010001;
12'b101111101001: finv2 = 23'b01010000100001100000010;
12'b101111101010: finv2 = 23'b01010000011011011110100;
12'b101111101011: finv2 = 23'b01010000010101011100111;
12'b101111101100: finv2 = 23'b01010000001111011011100;
12'b101111101101: finv2 = 23'b01010000001001011010001;
12'b101111101110: finv2 = 23'b01010000000011011001001;
12'b101111101111: finv2 = 23'b01001111111101011000001;
12'b101111110000: finv2 = 23'b01001111110111010111011;
12'b101111110001: finv2 = 23'b01001111110001010110110;
12'b101111110010: finv2 = 23'b01001111101011010110010;
12'b101111110011: finv2 = 23'b01001111100101010110000;
12'b101111110100: finv2 = 23'b01001111011111010101110;
12'b101111110101: finv2 = 23'b01001111011001010101111;
12'b101111110110: finv2 = 23'b01001111010011010110000;
12'b101111110111: finv2 = 23'b01001111001101010110011;
12'b101111111000: finv2 = 23'b01001111000111010110111;
12'b101111111001: finv2 = 23'b01001111000001010111100;
12'b101111111010: finv2 = 23'b01001110111011011000011;
12'b101111111011: finv2 = 23'b01001110110101011001011;
12'b101111111100: finv2 = 23'b01001110101111011010100;
12'b101111111101: finv2 = 23'b01001110101001011011110;
12'b101111111110: finv2 = 23'b01001110100011011101010;
12'b101111111111: finv2 = 23'b01001110011101011110111;
12'b110000000000: finv2 = 23'b01001110010111100000101;
12'b110000000001: finv2 = 23'b01001110010001100010101;
12'b110000000010: finv2 = 23'b01001110001011100100110;
12'b110000000011: finv2 = 23'b01001110000101100111000;
12'b110000000100: finv2 = 23'b01001101111111101001011;
12'b110000000101: finv2 = 23'b01001101111001101100000;
12'b110000000110: finv2 = 23'b01001101110011101110110;
12'b110000000111: finv2 = 23'b01001101101101110001101;
12'b110000001000: finv2 = 23'b01001101100111110100110;
12'b110000001001: finv2 = 23'b01001101100001110111111;
12'b110000001010: finv2 = 23'b01001101011011111011010;
12'b110000001011: finv2 = 23'b01001101010101111110111;
12'b110000001100: finv2 = 23'b01001101010000000010100;
12'b110000001101: finv2 = 23'b01001101001010000110011;
12'b110000001110: finv2 = 23'b01001101000100001010011;
12'b110000001111: finv2 = 23'b01001100111110001110101;
12'b110000010000: finv2 = 23'b01001100111000010010111;
12'b110000010001: finv2 = 23'b01001100110010010111011;
12'b110000010010: finv2 = 23'b01001100101100011100000;
12'b110000010011: finv2 = 23'b01001100100110100000111;
12'b110000010100: finv2 = 23'b01001100100000100101111;
12'b110000010101: finv2 = 23'b01001100011010101011000;
12'b110000010110: finv2 = 23'b01001100010100110000010;
12'b110000010111: finv2 = 23'b01001100001110110101110;
12'b110000011000: finv2 = 23'b01001100001000111011010;
12'b110000011001: finv2 = 23'b01001100000011000001000;
12'b110000011010: finv2 = 23'b01001011111101000111000;
12'b110000011011: finv2 = 23'b01001011110111001101000;
12'b110000011100: finv2 = 23'b01001011110001010011010;
12'b110000011101: finv2 = 23'b01001011101011011001101;
12'b110000011110: finv2 = 23'b01001011100101100000010;
12'b110000011111: finv2 = 23'b01001011011111100110111;
12'b110000100000: finv2 = 23'b01001011011001101101110;
12'b110000100001: finv2 = 23'b01001011010011110100110;
12'b110000100010: finv2 = 23'b01001011001101111100000;
12'b110000100011: finv2 = 23'b01001011001000000011010;
12'b110000100100: finv2 = 23'b01001011000010001010110;
12'b110000100101: finv2 = 23'b01001010111100010010011;
12'b110000100110: finv2 = 23'b01001010110110011010010;
12'b110000100111: finv2 = 23'b01001010110000100010001;
12'b110000101000: finv2 = 23'b01001010101010101010010;
12'b110000101001: finv2 = 23'b01001010100100110010100;
12'b110000101010: finv2 = 23'b01001010011110111011000;
12'b110000101011: finv2 = 23'b01001010011001000011101;
12'b110000101100: finv2 = 23'b01001010010011001100010;
12'b110000101101: finv2 = 23'b01001010001101010101010;
12'b110000101110: finv2 = 23'b01001010000111011110010;
12'b110000101111: finv2 = 23'b01001010000001100111100;
12'b110000110000: finv2 = 23'b01001001111011110000111;
12'b110000110001: finv2 = 23'b01001001110101111010011;
12'b110000110010: finv2 = 23'b01001001110000000100000;
12'b110000110011: finv2 = 23'b01001001101010001101111;
12'b110000110100: finv2 = 23'b01001001100100010111111;
12'b110000110101: finv2 = 23'b01001001011110100010000;
12'b110000110110: finv2 = 23'b01001001011000101100010;
12'b110000110111: finv2 = 23'b01001001010010110110110;
12'b110000111000: finv2 = 23'b01001001001101000001011;
12'b110000111001: finv2 = 23'b01001001000111001100001;
12'b110000111010: finv2 = 23'b01001001000001010111000;
12'b110000111011: finv2 = 23'b01001000111011100010001;
12'b110000111100: finv2 = 23'b01001000110101101101010;
12'b110000111101: finv2 = 23'b01001000101111111000110;
12'b110000111110: finv2 = 23'b01001000101010000100010;
12'b110000111111: finv2 = 23'b01001000100100001111111;
12'b110001000000: finv2 = 23'b01001000011110011011110;
12'b110001000001: finv2 = 23'b01001000011000100111110;
12'b110001000010: finv2 = 23'b01001000010010110011111;
12'b110001000011: finv2 = 23'b01001000001101000000010;
12'b110001000100: finv2 = 23'b01001000000111001100101;
12'b110001000101: finv2 = 23'b01001000000001011001010;
12'b110001000110: finv2 = 23'b01000111111011100110000;
12'b110001000111: finv2 = 23'b01000111110101110011000;
12'b110001001000: finv2 = 23'b01000111110000000000000;
12'b110001001001: finv2 = 23'b01000111101010001101010;
12'b110001001010: finv2 = 23'b01000111100100011010101;
12'b110001001011: finv2 = 23'b01000111011110101000010;
12'b110001001100: finv2 = 23'b01000111011000110101111;
12'b110001001101: finv2 = 23'b01000111010011000011110;
12'b110001001110: finv2 = 23'b01000111001101010001110;
12'b110001001111: finv2 = 23'b01000111000111011111111;
12'b110001010000: finv2 = 23'b01000111000001101110010;
12'b110001010001: finv2 = 23'b01000110111011111100101;
12'b110001010010: finv2 = 23'b01000110110110001011010;
12'b110001010011: finv2 = 23'b01000110110000011010000;
12'b110001010100: finv2 = 23'b01000110101010101001000;
12'b110001010101: finv2 = 23'b01000110100100111000000;
12'b110001010110: finv2 = 23'b01000110011111000111010;
12'b110001010111: finv2 = 23'b01000110011001010110101;
12'b110001011000: finv2 = 23'b01000110010011100110001;
12'b110001011001: finv2 = 23'b01000110001101110101110;
12'b110001011010: finv2 = 23'b01000110001000000101101;
12'b110001011011: finv2 = 23'b01000110000010010101101;
12'b110001011100: finv2 = 23'b01000101111100100101110;
12'b110001011101: finv2 = 23'b01000101110110110110000;
12'b110001011110: finv2 = 23'b01000101110001000110100;
12'b110001011111: finv2 = 23'b01000101101011010111001;
12'b110001100000: finv2 = 23'b01000101100101100111110;
12'b110001100001: finv2 = 23'b01000101011111111000110;
12'b110001100010: finv2 = 23'b01000101011010001001110;
12'b110001100011: finv2 = 23'b01000101010100011011000;
12'b110001100100: finv2 = 23'b01000101001110101100010;
12'b110001100101: finv2 = 23'b01000101001000111101110;
12'b110001100110: finv2 = 23'b01000101000011001111100;
12'b110001100111: finv2 = 23'b01000100111101100001010;
12'b110001101000: finv2 = 23'b01000100110111110011010;
12'b110001101001: finv2 = 23'b01000100110010000101010;
12'b110001101010: finv2 = 23'b01000100101100010111100;
12'b110001101011: finv2 = 23'b01000100100110101010000;
12'b110001101100: finv2 = 23'b01000100100000111100100;
12'b110001101101: finv2 = 23'b01000100011011001111010;
12'b110001101110: finv2 = 23'b01000100010101100010001;
12'b110001101111: finv2 = 23'b01000100001111110101001;
12'b110001110000: finv2 = 23'b01000100001010001000010;
12'b110001110001: finv2 = 23'b01000100000100011011100;
12'b110001110010: finv2 = 23'b01000011111110101111000;
12'b110001110011: finv2 = 23'b01000011111001000010101;
12'b110001110100: finv2 = 23'b01000011110011010110011;
12'b110001110101: finv2 = 23'b01000011101101101010010;
12'b110001110110: finv2 = 23'b01000011100111111110011;
12'b110001110111: finv2 = 23'b01000011100010010010100;
12'b110001111000: finv2 = 23'b01000011011100100110111;
12'b110001111001: finv2 = 23'b01000011010110111011011;
12'b110001111010: finv2 = 23'b01000011010001010000001;
12'b110001111011: finv2 = 23'b01000011001011100100111;
12'b110001111100: finv2 = 23'b01000011000101111001111;
12'b110001111101: finv2 = 23'b01000011000000001110111;
12'b110001111110: finv2 = 23'b01000010111010100100010;
12'b110001111111: finv2 = 23'b01000010110100111001101;
12'b110010000000: finv2 = 23'b01000010101111001111001;
12'b110010000001: finv2 = 23'b01000010101001100100111;
12'b110010000010: finv2 = 23'b01000010100011111010110;
12'b110010000011: finv2 = 23'b01000010011110010000110;
12'b110010000100: finv2 = 23'b01000010011000100110111;
12'b110010000101: finv2 = 23'b01000010010010111101001;
12'b110010000110: finv2 = 23'b01000010001101010011101;
12'b110010000111: finv2 = 23'b01000010000111101010001;
12'b110010001000: finv2 = 23'b01000010000010000000111;
12'b110010001001: finv2 = 23'b01000001111100010111111;
12'b110010001010: finv2 = 23'b01000001110110101110111;
12'b110010001011: finv2 = 23'b01000001110001000110000;
12'b110010001100: finv2 = 23'b01000001101011011101011;
12'b110010001101: finv2 = 23'b01000001100101110100111;
12'b110010001110: finv2 = 23'b01000001100000001100100;
12'b110010001111: finv2 = 23'b01000001011010100100010;
12'b110010010000: finv2 = 23'b01000001010100111100010;
12'b110010010001: finv2 = 23'b01000001001111010100010;
12'b110010010010: finv2 = 23'b01000001001001101100100;
12'b110010010011: finv2 = 23'b01000001000100000100111;
12'b110010010100: finv2 = 23'b01000000111110011101011;
12'b110010010101: finv2 = 23'b01000000111000110110000;
12'b110010010110: finv2 = 23'b01000000110011001110111;
12'b110010010111: finv2 = 23'b01000000101101100111111;
12'b110010011000: finv2 = 23'b01000000101000000000111;
12'b110010011001: finv2 = 23'b01000000100010011010001;
12'b110010011010: finv2 = 23'b01000000011100110011101;
12'b110010011011: finv2 = 23'b01000000010111001101001;
12'b110010011100: finv2 = 23'b01000000010001100110111;
12'b110010011101: finv2 = 23'b01000000001100000000101;
12'b110010011110: finv2 = 23'b01000000000110011010101;
12'b110010011111: finv2 = 23'b01000000000000110100110;
12'b110010100000: finv2 = 23'b00111111111011001111001;
12'b110010100001: finv2 = 23'b00111111110101101001100;
12'b110010100010: finv2 = 23'b00111111110000000100001;
12'b110010100011: finv2 = 23'b00111111101010011110110;
12'b110010100100: finv2 = 23'b00111111100100111001101;
12'b110010100101: finv2 = 23'b00111111011111010100101;
12'b110010100110: finv2 = 23'b00111111011001101111111;
12'b110010100111: finv2 = 23'b00111111010100001011001;
12'b110010101000: finv2 = 23'b00111111001110100110101;
12'b110010101001: finv2 = 23'b00111111001001000010001;
12'b110010101010: finv2 = 23'b00111111000011011101111;
12'b110010101011: finv2 = 23'b00111110111101111001110;
12'b110010101100: finv2 = 23'b00111110111000010101111;
12'b110010101101: finv2 = 23'b00111110110010110010000;
12'b110010101110: finv2 = 23'b00111110101101001110011;
12'b110010101111: finv2 = 23'b00111110100111101010110;
12'b110010110000: finv2 = 23'b00111110100010000111011;
12'b110010110001: finv2 = 23'b00111110011100100100001;
12'b110010110010: finv2 = 23'b00111110010111000001001;
12'b110010110011: finv2 = 23'b00111110010001011110001;
12'b110010110100: finv2 = 23'b00111110001011111011011;
12'b110010110101: finv2 = 23'b00111110000110011000101;
12'b110010110110: finv2 = 23'b00111110000000110110001;
12'b110010110111: finv2 = 23'b00111101111011010011110;
12'b110010111000: finv2 = 23'b00111101110101110001100;
12'b110010111001: finv2 = 23'b00111101110000001111100;
12'b110010111010: finv2 = 23'b00111101101010101101100;
12'b110010111011: finv2 = 23'b00111101100101001011110;
12'b110010111100: finv2 = 23'b00111101011111101010001;
12'b110010111101: finv2 = 23'b00111101011010001000101;
12'b110010111110: finv2 = 23'b00111101010100100111010;
12'b110010111111: finv2 = 23'b00111101001111000110000;
12'b110011000000: finv2 = 23'b00111101001001100100111;
12'b110011000001: finv2 = 23'b00111101000100000100000;
12'b110011000010: finv2 = 23'b00111100111110100011010;
12'b110011000011: finv2 = 23'b00111100111001000010101;
12'b110011000100: finv2 = 23'b00111100110011100010001;
12'b110011000101: finv2 = 23'b00111100101110000001110;
12'b110011000110: finv2 = 23'b00111100101000100001100;
12'b110011000111: finv2 = 23'b00111100100011000001100;
12'b110011001000: finv2 = 23'b00111100011101100001100;
12'b110011001001: finv2 = 23'b00111100011000000001110;
12'b110011001010: finv2 = 23'b00111100010010100010001;
12'b110011001011: finv2 = 23'b00111100001101000010101;
12'b110011001100: finv2 = 23'b00111100000111100011010;
12'b110011001101: finv2 = 23'b00111100000010000100000;
12'b110011001110: finv2 = 23'b00111011111100100101000;
12'b110011001111: finv2 = 23'b00111011110111000110000;
12'b110011010000: finv2 = 23'b00111011110001100111010;
12'b110011010001: finv2 = 23'b00111011101100001000101;
12'b110011010010: finv2 = 23'b00111011100110101010001;
12'b110011010011: finv2 = 23'b00111011100001001011110;
12'b110011010100: finv2 = 23'b00111011011011101101101;
12'b110011010101: finv2 = 23'b00111011010110001111100;
12'b110011010110: finv2 = 23'b00111011010000110001101;
12'b110011010111: finv2 = 23'b00111011001011010011110;
12'b110011011000: finv2 = 23'b00111011000101110110001;
12'b110011011001: finv2 = 23'b00111011000000011000101;
12'b110011011010: finv2 = 23'b00111010111010111011010;
12'b110011011011: finv2 = 23'b00111010110101011110001;
12'b110011011100: finv2 = 23'b00111010110000000001000;
12'b110011011101: finv2 = 23'b00111010101010100100001;
12'b110011011110: finv2 = 23'b00111010100101000111010;
12'b110011011111: finv2 = 23'b00111010011111101010101;
12'b110011100000: finv2 = 23'b00111010011010001110001;
12'b110011100001: finv2 = 23'b00111010010100110001110;
12'b110011100010: finv2 = 23'b00111010001111010101100;
12'b110011100011: finv2 = 23'b00111010001001111001100;
12'b110011100100: finv2 = 23'b00111010000100011101100;
12'b110011100101: finv2 = 23'b00111001111111000001110;
12'b110011100110: finv2 = 23'b00111001111001100110000;
12'b110011100111: finv2 = 23'b00111001110100001010100;
12'b110011101000: finv2 = 23'b00111001101110101111001;
12'b110011101001: finv2 = 23'b00111001101001010011111;
12'b110011101010: finv2 = 23'b00111001100011111000111;
12'b110011101011: finv2 = 23'b00111001011110011101111;
12'b110011101100: finv2 = 23'b00111001011001000011000;
12'b110011101101: finv2 = 23'b00111001010011101000011;
12'b110011101110: finv2 = 23'b00111001001110001101111;
12'b110011101111: finv2 = 23'b00111001001000110011100;
12'b110011110000: finv2 = 23'b00111001000011011001010;
12'b110011110001: finv2 = 23'b00111000111101111111001;
12'b110011110010: finv2 = 23'b00111000111000100101001;
12'b110011110011: finv2 = 23'b00111000110011001011010;
12'b110011110100: finv2 = 23'b00111000101101110001101;
12'b110011110101: finv2 = 23'b00111000101000011000000;
12'b110011110110: finv2 = 23'b00111000100010111110101;
12'b110011110111: finv2 = 23'b00111000011101100101011;
12'b110011111000: finv2 = 23'b00111000011000001100010;
12'b110011111001: finv2 = 23'b00111000010010110011010;
12'b110011111010: finv2 = 23'b00111000001101011010011;
12'b110011111011: finv2 = 23'b00111000001000000001101;
12'b110011111100: finv2 = 23'b00111000000010101001000;
12'b110011111101: finv2 = 23'b00110111111101010000101;
12'b110011111110: finv2 = 23'b00110111110111111000011;
12'b110011111111: finv2 = 23'b00110111110010100000001;
12'b110100000000: finv2 = 23'b00110111101101001000001;
12'b110100000001: finv2 = 23'b00110111100111110000010;
12'b110100000010: finv2 = 23'b00110111100010011000100;
12'b110100000011: finv2 = 23'b00110111011101000000111;
12'b110100000100: finv2 = 23'b00110111010111101001100;
12'b110100000101: finv2 = 23'b00110111010010010010001;
12'b110100000110: finv2 = 23'b00110111001100111011000;
12'b110100000111: finv2 = 23'b00110111000111100011111;
12'b110100001000: finv2 = 23'b00110111000010001101000;
12'b110100001001: finv2 = 23'b00110110111100110110010;
12'b110100001010: finv2 = 23'b00110110110111011111101;
12'b110100001011: finv2 = 23'b00110110110010001001001;
12'b110100001100: finv2 = 23'b00110110101100110010110;
12'b110100001101: finv2 = 23'b00110110100111011100100;
12'b110100001110: finv2 = 23'b00110110100010000110011;
12'b110100001111: finv2 = 23'b00110110011100110000100;
12'b110100010000: finv2 = 23'b00110110010111011010101;
12'b110100010001: finv2 = 23'b00110110010010000101000;
12'b110100010010: finv2 = 23'b00110110001100101111100;
12'b110100010011: finv2 = 23'b00110110000111011010001;
12'b110100010100: finv2 = 23'b00110110000010000100111;
12'b110100010101: finv2 = 23'b00110101111100101111110;
12'b110100010110: finv2 = 23'b00110101110111011010110;
12'b110100010111: finv2 = 23'b00110101110010000101111;
12'b110100011000: finv2 = 23'b00110101101100110001010;
12'b110100011001: finv2 = 23'b00110101100111011100101;
12'b110100011010: finv2 = 23'b00110101100010001000010;
12'b110100011011: finv2 = 23'b00110101011100110011111;
12'b110100011100: finv2 = 23'b00110101010111011111110;
12'b110100011101: finv2 = 23'b00110101010010001011110;
12'b110100011110: finv2 = 23'b00110101001100110111111;
12'b110100011111: finv2 = 23'b00110101000111100100001;
12'b110100100000: finv2 = 23'b00110101000010010000100;
12'b110100100001: finv2 = 23'b00110100111100111101000;
12'b110100100010: finv2 = 23'b00110100110111101001101;
12'b110100100011: finv2 = 23'b00110100110010010110100;
12'b110100100100: finv2 = 23'b00110100101101000011011;
12'b110100100101: finv2 = 23'b00110100100111110000100;
12'b110100100110: finv2 = 23'b00110100100010011101110;
12'b110100100111: finv2 = 23'b00110100011101001011000;
12'b110100101000: finv2 = 23'b00110100010111111000100;
12'b110100101001: finv2 = 23'b00110100010010100110001;
12'b110100101010: finv2 = 23'b00110100001101010011111;
12'b110100101011: finv2 = 23'b00110100001000000001110;
12'b110100101100: finv2 = 23'b00110100000010101111110;
12'b110100101101: finv2 = 23'b00110011111101011110000;
12'b110100101110: finv2 = 23'b00110011111000001100010;
12'b110100101111: finv2 = 23'b00110011110010111010110;
12'b110100110000: finv2 = 23'b00110011101101101001010;
12'b110100110001: finv2 = 23'b00110011101000011000000;
12'b110100110010: finv2 = 23'b00110011100011000110110;
12'b110100110011: finv2 = 23'b00110011011101110101110;
12'b110100110100: finv2 = 23'b00110011011000100100111;
12'b110100110101: finv2 = 23'b00110011010011010100001;
12'b110100110110: finv2 = 23'b00110011001110000011100;
12'b110100110111: finv2 = 23'b00110011001000110011000;
12'b110100111000: finv2 = 23'b00110011000011100010101;
12'b110100111001: finv2 = 23'b00110010111110010010100;
12'b110100111010: finv2 = 23'b00110010111001000010011;
12'b110100111011: finv2 = 23'b00110010110011110010011;
12'b110100111100: finv2 = 23'b00110010101110100010101;
12'b110100111101: finv2 = 23'b00110010101001010011000;
12'b110100111110: finv2 = 23'b00110010100100000011011;
12'b110100111111: finv2 = 23'b00110010011110110100000;
12'b110101000000: finv2 = 23'b00110010011001100100110;
12'b110101000001: finv2 = 23'b00110010010100010101101;
12'b110101000010: finv2 = 23'b00110010001111000110101;
12'b110101000011: finv2 = 23'b00110010001001110111110;
12'b110101000100: finv2 = 23'b00110010000100101001000;
12'b110101000101: finv2 = 23'b00110001111111011010011;
12'b110101000110: finv2 = 23'b00110001111010001011111;
12'b110101000111: finv2 = 23'b00110001110100111101101;
12'b110101001000: finv2 = 23'b00110001101111101111011;
12'b110101001001: finv2 = 23'b00110001101010100001010;
12'b110101001010: finv2 = 23'b00110001100101010011011;
12'b110101001011: finv2 = 23'b00110001100000000101101;
12'b110101001100: finv2 = 23'b00110001011010110111111;
12'b110101001101: finv2 = 23'b00110001010101101010011;
12'b110101001110: finv2 = 23'b00110001010000011101000;
12'b110101001111: finv2 = 23'b00110001001011001111110;
12'b110101010000: finv2 = 23'b00110001000110000010101;
12'b110101010001: finv2 = 23'b00110001000000110101101;
12'b110101010010: finv2 = 23'b00110000111011101000110;
12'b110101010011: finv2 = 23'b00110000110110011100000;
12'b110101010100: finv2 = 23'b00110000110001001111011;
12'b110101010101: finv2 = 23'b00110000101100000010111;
12'b110101010110: finv2 = 23'b00110000100110110110100;
12'b110101010111: finv2 = 23'b00110000100001101010011;
12'b110101011000: finv2 = 23'b00110000011100011110010;
12'b110101011001: finv2 = 23'b00110000010111010010011;
12'b110101011010: finv2 = 23'b00110000010010000110100;
12'b110101011011: finv2 = 23'b00110000001100111010111;
12'b110101011100: finv2 = 23'b00110000000111101111011;
12'b110101011101: finv2 = 23'b00110000000010100011111;
12'b110101011110: finv2 = 23'b00101111111101011000101;
12'b110101011111: finv2 = 23'b00101111111000001101100;
12'b110101100000: finv2 = 23'b00101111110011000010100;
12'b110101100001: finv2 = 23'b00101111101101110111101;
12'b110101100010: finv2 = 23'b00101111101000101100111;
12'b110101100011: finv2 = 23'b00101111100011100010010;
12'b110101100100: finv2 = 23'b00101111011110010111110;
12'b110101100101: finv2 = 23'b00101111011001001101011;
12'b110101100110: finv2 = 23'b00101111010100000011010;
12'b110101100111: finv2 = 23'b00101111001110111001001;
12'b110101101000: finv2 = 23'b00101111001001101111001;
12'b110101101001: finv2 = 23'b00101111000100100101011;
12'b110101101010: finv2 = 23'b00101110111111011011101;
12'b110101101011: finv2 = 23'b00101110111010010010001;
12'b110101101100: finv2 = 23'b00101110110101001000101;
12'b110101101101: finv2 = 23'b00101110101111111111011;
12'b110101101110: finv2 = 23'b00101110101010110110001;
12'b110101101111: finv2 = 23'b00101110100101101101001;
12'b110101110000: finv2 = 23'b00101110100000100100010;
12'b110101110001: finv2 = 23'b00101110011011011011100;
12'b110101110010: finv2 = 23'b00101110010110010010110;
12'b110101110011: finv2 = 23'b00101110010001001010010;
12'b110101110100: finv2 = 23'b00101110001100000001111;
12'b110101110101: finv2 = 23'b00101110000110111001101;
12'b110101110110: finv2 = 23'b00101110000001110001100;
12'b110101110111: finv2 = 23'b00101101111100101001100;
12'b110101111000: finv2 = 23'b00101101110111100001101;
12'b110101111001: finv2 = 23'b00101101110010011001111;
12'b110101111010: finv2 = 23'b00101101101101010010011;
12'b110101111011: finv2 = 23'b00101101101000001010111;
12'b110101111100: finv2 = 23'b00101101100011000011100;
12'b110101111101: finv2 = 23'b00101101011101111100010;
12'b110101111110: finv2 = 23'b00101101011000110101010;
12'b110101111111: finv2 = 23'b00101101010011101110010;
12'b110110000000: finv2 = 23'b00101101001110100111100;
12'b110110000001: finv2 = 23'b00101101001001100000110;
12'b110110000010: finv2 = 23'b00101101000100011010010;
12'b110110000011: finv2 = 23'b00101100111111010011110;
12'b110110000100: finv2 = 23'b00101100111010001101100;
12'b110110000101: finv2 = 23'b00101100110101000111010;
12'b110110000110: finv2 = 23'b00101100110000000001010;
12'b110110000111: finv2 = 23'b00101100101010111011011;
12'b110110001000: finv2 = 23'b00101100100101110101100;
12'b110110001001: finv2 = 23'b00101100100000101111111;
12'b110110001010: finv2 = 23'b00101100011011101010011;
12'b110110001011: finv2 = 23'b00101100010110100101000;
12'b110110001100: finv2 = 23'b00101100010001011111110;
12'b110110001101: finv2 = 23'b00101100001100011010101;
12'b110110001110: finv2 = 23'b00101100000111010101100;
12'b110110001111: finv2 = 23'b00101100000010010000101;
12'b110110010000: finv2 = 23'b00101011111101001011111;
12'b110110010001: finv2 = 23'b00101011111000000111010;
12'b110110010010: finv2 = 23'b00101011110011000010110;
12'b110110010011: finv2 = 23'b00101011101101111110100;
12'b110110010100: finv2 = 23'b00101011101000111010010;
12'b110110010101: finv2 = 23'b00101011100011110110001;
12'b110110010110: finv2 = 23'b00101011011110110010001;
12'b110110010111: finv2 = 23'b00101011011001101110010;
12'b110110011000: finv2 = 23'b00101011010100101010100;
12'b110110011001: finv2 = 23'b00101011001111100110111;
12'b110110011010: finv2 = 23'b00101011001010100011100;
12'b110110011011: finv2 = 23'b00101011000101100000001;
12'b110110011100: finv2 = 23'b00101011000000011100111;
12'b110110011101: finv2 = 23'b00101010111011011001111;
12'b110110011110: finv2 = 23'b00101010110110010110111;
12'b110110011111: finv2 = 23'b00101010110001010100000;
12'b110110100000: finv2 = 23'b00101010101100010001011;
12'b110110100001: finv2 = 23'b00101010100111001110110;
12'b110110100010: finv2 = 23'b00101010100010001100011;
12'b110110100011: finv2 = 23'b00101010011101001010000;
12'b110110100100: finv2 = 23'b00101010011000000111110;
12'b110110100101: finv2 = 23'b00101010010011000101110;
12'b110110100110: finv2 = 23'b00101010001110000011110;
12'b110110100111: finv2 = 23'b00101010001001000010000;
12'b110110101000: finv2 = 23'b00101010000100000000011;
12'b110110101001: finv2 = 23'b00101001111110111110110;
12'b110110101010: finv2 = 23'b00101001111001111101011;
12'b110110101011: finv2 = 23'b00101001110100111100000;
12'b110110101100: finv2 = 23'b00101001101111111010111;
12'b110110101101: finv2 = 23'b00101001101010111001111;
12'b110110101110: finv2 = 23'b00101001100101111000111;
12'b110110101111: finv2 = 23'b00101001100000111000001;
12'b110110110000: finv2 = 23'b00101001011011110111011;
12'b110110110001: finv2 = 23'b00101001010110110110111;
12'b110110110010: finv2 = 23'b00101001010001110110100;
12'b110110110011: finv2 = 23'b00101001001100110110010;
12'b110110110100: finv2 = 23'b00101001000111110110000;
12'b110110110101: finv2 = 23'b00101001000010110110000;
12'b110110110110: finv2 = 23'b00101000111101110110001;
12'b110110110111: finv2 = 23'b00101000111000110110010;
12'b110110111000: finv2 = 23'b00101000110011110110101;
12'b110110111001: finv2 = 23'b00101000101110110111001;
12'b110110111010: finv2 = 23'b00101000101001110111110;
12'b110110111011: finv2 = 23'b00101000100100111000011;
12'b110110111100: finv2 = 23'b00101000011111111001010;
12'b110110111101: finv2 = 23'b00101000011010111010010;
12'b110110111110: finv2 = 23'b00101000010101111011011;
12'b110110111111: finv2 = 23'b00101000010000111100101;
12'b110111000000: finv2 = 23'b00101000001011111101111;
12'b110111000001: finv2 = 23'b00101000000110111111011;
12'b110111000010: finv2 = 23'b00101000000010000001000;
12'b110111000011: finv2 = 23'b00100111111101000010110;
12'b110111000100: finv2 = 23'b00100111111000000100101;
12'b110111000101: finv2 = 23'b00100111110011000110100;
12'b110111000110: finv2 = 23'b00100111101110001000101;
12'b110111000111: finv2 = 23'b00100111101001001010111;
12'b110111001000: finv2 = 23'b00100111100100001101010;
12'b110111001001: finv2 = 23'b00100111011111001111110;
12'b110111001010: finv2 = 23'b00100111011010010010010;
12'b110111001011: finv2 = 23'b00100111010101010101000;
12'b110111001100: finv2 = 23'b00100111010000010111111;
12'b110111001101: finv2 = 23'b00100111001011011010111;
12'b110111001110: finv2 = 23'b00100111000110011110000;
12'b110111001111: finv2 = 23'b00100111000001100001001;
12'b110111010000: finv2 = 23'b00100110111100100100100;
12'b110111010001: finv2 = 23'b00100110110111101000000;
12'b110111010010: finv2 = 23'b00100110110010101011101;
12'b110111010011: finv2 = 23'b00100110101101101111011;
12'b110111010100: finv2 = 23'b00100110101000110011001;
12'b110111010101: finv2 = 23'b00100110100011110111001;
12'b110111010110: finv2 = 23'b00100110011110111011010;
12'b110111010111: finv2 = 23'b00100110011001111111100;
12'b110111011000: finv2 = 23'b00100110010101000011110;
12'b110111011001: finv2 = 23'b00100110010000001000010;
12'b110111011010: finv2 = 23'b00100110001011001100111;
12'b110111011011: finv2 = 23'b00100110000110010001101;
12'b110111011100: finv2 = 23'b00100110000001010110011;
12'b110111011101: finv2 = 23'b00100101111100011011011;
12'b110111011110: finv2 = 23'b00100101110111100000100;
12'b110111011111: finv2 = 23'b00100101110010100101101;
12'b110111100000: finv2 = 23'b00100101101101101011000;
12'b110111100001: finv2 = 23'b00100101101000110000100;
12'b110111100010: finv2 = 23'b00100101100011110110000;
12'b110111100011: finv2 = 23'b00100101011110111011110;
12'b110111100100: finv2 = 23'b00100101011010000001101;
12'b110111100101: finv2 = 23'b00100101010101000111100;
12'b110111100110: finv2 = 23'b00100101010000001101101;
12'b110111100111: finv2 = 23'b00100101001011010011110;
12'b110111101000: finv2 = 23'b00100101000110011010001;
12'b110111101001: finv2 = 23'b00100101000001100000100;
12'b110111101010: finv2 = 23'b00100100111100100111001;
12'b110111101011: finv2 = 23'b00100100110111101101110;
12'b110111101100: finv2 = 23'b00100100110010110100101;
12'b110111101101: finv2 = 23'b00100100101101111011100;
12'b110111101110: finv2 = 23'b00100100101001000010101;
12'b110111101111: finv2 = 23'b00100100100100001001110;
12'b110111110000: finv2 = 23'b00100100011111010001001;
12'b110111110001: finv2 = 23'b00100100011010011000100;
12'b110111110010: finv2 = 23'b00100100010101100000000;
12'b110111110011: finv2 = 23'b00100100010000100111110;
12'b110111110100: finv2 = 23'b00100100001011101111100;
12'b110111110101: finv2 = 23'b00100100000110110111011;
12'b110111110110: finv2 = 23'b00100100000001111111100;
12'b110111110111: finv2 = 23'b00100011111101000111101;
12'b110111111000: finv2 = 23'b00100011111000001111111;
12'b110111111001: finv2 = 23'b00100011110011011000010;
12'b110111111010: finv2 = 23'b00100011101110100000110;
12'b110111111011: finv2 = 23'b00100011101001101001011;
12'b110111111100: finv2 = 23'b00100011100100110010010;
12'b110111111101: finv2 = 23'b00100011011111111011001;
12'b110111111110: finv2 = 23'b00100011011011000100001;
12'b110111111111: finv2 = 23'b00100011010110001101010;
12'b111000000000: finv2 = 23'b00100011010001010110100;
12'b111000000001: finv2 = 23'b00100011001100011111111;
12'b111000000010: finv2 = 23'b00100011000111101001011;
12'b111000000011: finv2 = 23'b00100011000010110011000;
12'b111000000100: finv2 = 23'b00100010111101111100101;
12'b111000000101: finv2 = 23'b00100010111001000110100;
12'b111000000110: finv2 = 23'b00100010110100010000100;
12'b111000000111: finv2 = 23'b00100010101111011010101;
12'b111000001000: finv2 = 23'b00100010101010100100111;
12'b111000001001: finv2 = 23'b00100010100101101111001;
12'b111000001010: finv2 = 23'b00100010100000111001101;
12'b111000001011: finv2 = 23'b00100010011100000100010;
12'b111000001100: finv2 = 23'b00100010010111001110111;
12'b111000001101: finv2 = 23'b00100010010010011001110;
12'b111000001110: finv2 = 23'b00100010001101100100101;
12'b111000001111: finv2 = 23'b00100010001000101111110;
12'b111000010000: finv2 = 23'b00100010000011111010111;
12'b111000010001: finv2 = 23'b00100001111111000110010;
12'b111000010010: finv2 = 23'b00100001111010010001101;
12'b111000010011: finv2 = 23'b00100001110101011101010;
12'b111000010100: finv2 = 23'b00100001110000101000111;
12'b111000010101: finv2 = 23'b00100001101011110100101;
12'b111000010110: finv2 = 23'b00100001100111000000101;
12'b111000010111: finv2 = 23'b00100001100010001100101;
12'b111000011000: finv2 = 23'b00100001011101011000110;
12'b111000011001: finv2 = 23'b00100001011000100101000;
12'b111000011010: finv2 = 23'b00100001010011110001011;
12'b111000011011: finv2 = 23'b00100001001110111101111;
12'b111000011100: finv2 = 23'b00100001001010001010100;
12'b111000011101: finv2 = 23'b00100001000101010111010;
12'b111000011110: finv2 = 23'b00100001000000100100001;
12'b111000011111: finv2 = 23'b00100000111011110001001;
12'b111000100000: finv2 = 23'b00100000110110111110010;
12'b111000100001: finv2 = 23'b00100000110010001011011;
12'b111000100010: finv2 = 23'b00100000101101011000110;
12'b111000100011: finv2 = 23'b00100000101000100110010;
12'b111000100100: finv2 = 23'b00100000100011110011111;
12'b111000100101: finv2 = 23'b00100000011111000001100;
12'b111000100110: finv2 = 23'b00100000011010001111011;
12'b111000100111: finv2 = 23'b00100000010101011101010;
12'b111000101000: finv2 = 23'b00100000010000101011011;
12'b111000101001: finv2 = 23'b00100000001011111001100;
12'b111000101010: finv2 = 23'b00100000000111000111110;
12'b111000101011: finv2 = 23'b00100000000010010110010;
12'b111000101100: finv2 = 23'b00011111111101100100110;
12'b111000101101: finv2 = 23'b00011111111000110011011;
12'b111000101110: finv2 = 23'b00011111110100000010001;
12'b111000101111: finv2 = 23'b00011111101111010001000;
12'b111000110000: finv2 = 23'b00011111101010100000000;
12'b111000110001: finv2 = 23'b00011111100101101111001;
12'b111000110010: finv2 = 23'b00011111100000111110011;
12'b111000110011: finv2 = 23'b00011111011100001101110;
12'b111000110100: finv2 = 23'b00011111010111011101010;
12'b111000110101: finv2 = 23'b00011111010010101100111;
12'b111000110110: finv2 = 23'b00011111001101111100100;
12'b111000110111: finv2 = 23'b00011111001001001100011;
12'b111000111000: finv2 = 23'b00011111000100011100011;
12'b111000111001: finv2 = 23'b00011110111111101100011;
12'b111000111010: finv2 = 23'b00011110111010111100101;
12'b111000111011: finv2 = 23'b00011110110110001100111;
12'b111000111100: finv2 = 23'b00011110110001011101011;
12'b111000111101: finv2 = 23'b00011110101100101101111;
12'b111000111110: finv2 = 23'b00011110100111111110100;
12'b111000111111: finv2 = 23'b00011110100011001111010;
12'b111001000000: finv2 = 23'b00011110011110100000001;
12'b111001000001: finv2 = 23'b00011110011001110001010;
12'b111001000010: finv2 = 23'b00011110010101000010011;
12'b111001000011: finv2 = 23'b00011110010000010011100;
12'b111001000100: finv2 = 23'b00011110001011100100111;
12'b111001000101: finv2 = 23'b00011110000110110110011;
12'b111001000110: finv2 = 23'b00011110000010001000000;
12'b111001000111: finv2 = 23'b00011101111101011001110;
12'b111001001000: finv2 = 23'b00011101111000101011100;
12'b111001001001: finv2 = 23'b00011101110011111101100;
12'b111001001010: finv2 = 23'b00011101101111001111100;
12'b111001001011: finv2 = 23'b00011101101010100001110;
12'b111001001100: finv2 = 23'b00011101100101110100000;
12'b111001001101: finv2 = 23'b00011101100001000110011;
12'b111001001110: finv2 = 23'b00011101011100011001000;
12'b111001001111: finv2 = 23'b00011101010111101011101;
12'b111001010000: finv2 = 23'b00011101010010111110011;
12'b111001010001: finv2 = 23'b00011101001110010001010;
12'b111001010010: finv2 = 23'b00011101001001100100010;
12'b111001010011: finv2 = 23'b00011101000100110111011;
12'b111001010100: finv2 = 23'b00011101000000001010101;
12'b111001010101: finv2 = 23'b00011100111011011101111;
12'b111001010110: finv2 = 23'b00011100110110110001011;
12'b111001010111: finv2 = 23'b00011100110010000101000;
12'b111001011000: finv2 = 23'b00011100101101011000101;
12'b111001011001: finv2 = 23'b00011100101000101100100;
12'b111001011010: finv2 = 23'b00011100100100000000011;
12'b111001011011: finv2 = 23'b00011100011111010100011;
12'b111001011100: finv2 = 23'b00011100011010101000101;
12'b111001011101: finv2 = 23'b00011100010101111100111;
12'b111001011110: finv2 = 23'b00011100010001010001010;
12'b111001011111: finv2 = 23'b00011100001100100101110;
12'b111001100000: finv2 = 23'b00011100000111111010011;
12'b111001100001: finv2 = 23'b00011100000011001111001;
12'b111001100010: finv2 = 23'b00011011111110100100000;
12'b111001100011: finv2 = 23'b00011011111001111000111;
12'b111001100100: finv2 = 23'b00011011110101001110000;
12'b111001100101: finv2 = 23'b00011011110000100011010;
12'b111001100110: finv2 = 23'b00011011101011111000100;
12'b111001100111: finv2 = 23'b00011011100111001101111;
12'b111001101000: finv2 = 23'b00011011100010100011100;
12'b111001101001: finv2 = 23'b00011011011101111001001;
12'b111001101010: finv2 = 23'b00011011011001001110111;
12'b111001101011: finv2 = 23'b00011011010100100100110;
12'b111001101100: finv2 = 23'b00011011001111111010110;
12'b111001101101: finv2 = 23'b00011011001011010000111;
12'b111001101110: finv2 = 23'b00011011000110100111001;
12'b111001101111: finv2 = 23'b00011011000001111101100;
12'b111001110000: finv2 = 23'b00011010111101010011111;
12'b111001110001: finv2 = 23'b00011010111000101010100;
12'b111001110010: finv2 = 23'b00011010110100000001010;
12'b111001110011: finv2 = 23'b00011010101111011000000;
12'b111001110100: finv2 = 23'b00011010101010101110111;
12'b111001110101: finv2 = 23'b00011010100110000110000;
12'b111001110110: finv2 = 23'b00011010100001011101001;
12'b111001110111: finv2 = 23'b00011010011100110100011;
12'b111001111000: finv2 = 23'b00011010011000001011110;
12'b111001111001: finv2 = 23'b00011010010011100011010;
12'b111001111010: finv2 = 23'b00011010001110111010111;
12'b111001111011: finv2 = 23'b00011010001010010010100;
12'b111001111100: finv2 = 23'b00011010000101101010011;
12'b111001111101: finv2 = 23'b00011010000001000010010;
12'b111001111110: finv2 = 23'b00011001111100011010011;
12'b111001111111: finv2 = 23'b00011001110111110010100;
12'b111010000000: finv2 = 23'b00011001110011001010111;
12'b111010000001: finv2 = 23'b00011001101110100011010;
12'b111010000010: finv2 = 23'b00011001101001111011110;
12'b111010000011: finv2 = 23'b00011001100101010100011;
12'b111010000100: finv2 = 23'b00011001100000101101001;
12'b111010000101: finv2 = 23'b00011001011100000110000;
12'b111010000110: finv2 = 23'b00011001010111011110111;
12'b111010000111: finv2 = 23'b00011001010010111000000;
12'b111010001000: finv2 = 23'b00011001001110010001001;
12'b111010001001: finv2 = 23'b00011001001001101010100;
12'b111010001010: finv2 = 23'b00011001000101000011111;
12'b111010001011: finv2 = 23'b00011001000000011101011;
12'b111010001100: finv2 = 23'b00011000111011110111001;
12'b111010001101: finv2 = 23'b00011000110111010000111;
12'b111010001110: finv2 = 23'b00011000110010101010110;
12'b111010001111: finv2 = 23'b00011000101110000100110;
12'b111010010000: finv2 = 23'b00011000101001011110110;
12'b111010010001: finv2 = 23'b00011000100100111001000;
12'b111010010010: finv2 = 23'b00011000100000010011010;
12'b111010010011: finv2 = 23'b00011000011011101101110;
12'b111010010100: finv2 = 23'b00011000010111001000010;
12'b111010010101: finv2 = 23'b00011000010010100011000;
12'b111010010110: finv2 = 23'b00011000001101111101110;
12'b111010010111: finv2 = 23'b00011000001001011000101;
12'b111010011000: finv2 = 23'b00011000000100110011101;
12'b111010011001: finv2 = 23'b00011000000000001110110;
12'b111010011010: finv2 = 23'b00010111111011101001111;
12'b111010011011: finv2 = 23'b00010111110111000101010;
12'b111010011100: finv2 = 23'b00010111110010100000110;
12'b111010011101: finv2 = 23'b00010111101101111100010;
12'b111010011110: finv2 = 23'b00010111101001010111111;
12'b111010011111: finv2 = 23'b00010111100100110011110;
12'b111010100000: finv2 = 23'b00010111100000001111101;
12'b111010100001: finv2 = 23'b00010111011011101011101;
12'b111010100010: finv2 = 23'b00010111010111000111110;
12'b111010100011: finv2 = 23'b00010111010010100011111;
12'b111010100100: finv2 = 23'b00010111001110000000010;
12'b111010100101: finv2 = 23'b00010111001001011100110;
12'b111010100110: finv2 = 23'b00010111000100111001010;
12'b111010100111: finv2 = 23'b00010111000000010110000;
12'b111010101000: finv2 = 23'b00010110111011110010110;
12'b111010101001: finv2 = 23'b00010110110111001111101;
12'b111010101010: finv2 = 23'b00010110110010101100101;
12'b111010101011: finv2 = 23'b00010110101110001001110;
12'b111010101100: finv2 = 23'b00010110101001100111000;
12'b111010101101: finv2 = 23'b00010110100101000100011;
12'b111010101110: finv2 = 23'b00010110100000100001110;
12'b111010101111: finv2 = 23'b00010110011011111111011;
12'b111010110000: finv2 = 23'b00010110010111011101000;
12'b111010110001: finv2 = 23'b00010110010010111010110;
12'b111010110010: finv2 = 23'b00010110001110011000110;
12'b111010110011: finv2 = 23'b00010110001001110110110;
12'b111010110100: finv2 = 23'b00010110000101010100110;
12'b111010110101: finv2 = 23'b00010110000000110011000;
12'b111010110110: finv2 = 23'b00010101111100010001011;
12'b111010110111: finv2 = 23'b00010101110111101111111;
12'b111010111000: finv2 = 23'b00010101110011001110011;
12'b111010111001: finv2 = 23'b00010101101110101101000;
12'b111010111010: finv2 = 23'b00010101101010001011111;
12'b111010111011: finv2 = 23'b00010101100101101010110;
12'b111010111100: finv2 = 23'b00010101100001001001110;
12'b111010111101: finv2 = 23'b00010101011100101000111;
12'b111010111110: finv2 = 23'b00010101011000001000000;
12'b111010111111: finv2 = 23'b00010101010011100111011;
12'b111011000000: finv2 = 23'b00010101001111000110110;
12'b111011000001: finv2 = 23'b00010101001010100110011;
12'b111011000010: finv2 = 23'b00010101000110000110000;
12'b111011000011: finv2 = 23'b00010101000001100101110;
12'b111011000100: finv2 = 23'b00010100111101000101101;
12'b111011000101: finv2 = 23'b00010100111000100101101;
12'b111011000110: finv2 = 23'b00010100110100000101110;
12'b111011000111: finv2 = 23'b00010100101111100110000;
12'b111011001000: finv2 = 23'b00010100101011000110010;
12'b111011001001: finv2 = 23'b00010100100110100110110;
12'b111011001010: finv2 = 23'b00010100100010000111010;
12'b111011001011: finv2 = 23'b00010100011101100111111;
12'b111011001100: finv2 = 23'b00010100011001001000101;
12'b111011001101: finv2 = 23'b00010100010100101001100;
12'b111011001110: finv2 = 23'b00010100010000001010100;
12'b111011001111: finv2 = 23'b00010100001011101011100;
12'b111011010000: finv2 = 23'b00010100000111001100110;
12'b111011010001: finv2 = 23'b00010100000010101110000;
12'b111011010010: finv2 = 23'b00010011111110001111100;
12'b111011010011: finv2 = 23'b00010011111001110001000;
12'b111011010100: finv2 = 23'b00010011110101010010101;
12'b111011010101: finv2 = 23'b00010011110000110100011;
12'b111011010110: finv2 = 23'b00010011101100010110010;
12'b111011010111: finv2 = 23'b00010011100111111000001;
12'b111011011000: finv2 = 23'b00010011100011011010010;
12'b111011011001: finv2 = 23'b00010011011110111100011;
12'b111011011010: finv2 = 23'b00010011011010011110101;
12'b111011011011: finv2 = 23'b00010011010110000001000;
12'b111011011100: finv2 = 23'b00010011010001100011100;
12'b111011011101: finv2 = 23'b00010011001101000110001;
12'b111011011110: finv2 = 23'b00010011001000101000111;
12'b111011011111: finv2 = 23'b00010011000100001011101;
12'b111011100000: finv2 = 23'b00010010111111101110101;
12'b111011100001: finv2 = 23'b00010010111011010001101;
12'b111011100010: finv2 = 23'b00010010110110110100110;
12'b111011100011: finv2 = 23'b00010010110010011000000;
12'b111011100100: finv2 = 23'b00010010101101111011011;
12'b111011100101: finv2 = 23'b00010010101001011110111;
12'b111011100110: finv2 = 23'b00010010100101000010100;
12'b111011100111: finv2 = 23'b00010010100000100110001;
12'b111011101000: finv2 = 23'b00010010011100001010000;
12'b111011101001: finv2 = 23'b00010010010111101101111;
12'b111011101010: finv2 = 23'b00010010010011010001111;
12'b111011101011: finv2 = 23'b00010010001110110110000;
12'b111011101100: finv2 = 23'b00010010001010011010010;
12'b111011101101: finv2 = 23'b00010010000101111110100;
12'b111011101110: finv2 = 23'b00010010000001100011000;
12'b111011101111: finv2 = 23'b00010001111101000111100;
12'b111011110000: finv2 = 23'b00010001111000101100001;
12'b111011110001: finv2 = 23'b00010001110100010000111;
12'b111011110010: finv2 = 23'b00010001101111110101110;
12'b111011110011: finv2 = 23'b00010001101011011010110;
12'b111011110100: finv2 = 23'b00010001100110111111111;
12'b111011110101: finv2 = 23'b00010001100010100101000;
12'b111011110110: finv2 = 23'b00010001011110001010011;
12'b111011110111: finv2 = 23'b00010001011001101111110;
12'b111011111000: finv2 = 23'b00010001010101010101010;
12'b111011111001: finv2 = 23'b00010001010000111010111;
12'b111011111010: finv2 = 23'b00010001001100100000101;
12'b111011111011: finv2 = 23'b00010001001000000110011;
12'b111011111100: finv2 = 23'b00010001000011101100011;
12'b111011111101: finv2 = 23'b00010000111111010010011;
12'b111011111110: finv2 = 23'b00010000111010111000101;
12'b111011111111: finv2 = 23'b00010000110110011110111;
12'b111100000000: finv2 = 23'b00010000110010000101010;
12'b111100000001: finv2 = 23'b00010000101101101011101;
12'b111100000010: finv2 = 23'b00010000101001010010010;
12'b111100000011: finv2 = 23'b00010000100100111000111;
12'b111100000100: finv2 = 23'b00010000100000011111110;
12'b111100000101: finv2 = 23'b00010000011100000110101;
12'b111100000110: finv2 = 23'b00010000010111101101101;
12'b111100000111: finv2 = 23'b00010000010011010100110;
12'b111100001000: finv2 = 23'b00010000001110111100000;
12'b111100001001: finv2 = 23'b00010000001010100011010;
12'b111100001010: finv2 = 23'b00010000000110001010110;
12'b111100001011: finv2 = 23'b00010000000001110010010;
12'b111100001100: finv2 = 23'b00001111111101011001111;
12'b111100001101: finv2 = 23'b00001111111001000001101;
12'b111100001110: finv2 = 23'b00001111110100101001100;
12'b111100001111: finv2 = 23'b00001111110000010001011;
12'b111100010000: finv2 = 23'b00001111101011111001100;
12'b111100010001: finv2 = 23'b00001111100111100001101;
12'b111100010010: finv2 = 23'b00001111100011001001111;
12'b111100010011: finv2 = 23'b00001111011110110010010;
12'b111100010100: finv2 = 23'b00001111011010011010110;
12'b111100010101: finv2 = 23'b00001111010110000011011;
12'b111100010110: finv2 = 23'b00001111010001101100000;
12'b111100010111: finv2 = 23'b00001111001101010100111;
12'b111100011000: finv2 = 23'b00001111001000111101110;
12'b111100011001: finv2 = 23'b00001111000100100110110;
12'b111100011010: finv2 = 23'b00001111000000001111111;
12'b111100011011: finv2 = 23'b00001110111011111001001;
12'b111100011100: finv2 = 23'b00001110110111100010011;
12'b111100011101: finv2 = 23'b00001110110011001011111;
12'b111100011110: finv2 = 23'b00001110101110110101011;
12'b111100011111: finv2 = 23'b00001110101010011111000;
12'b111100100000: finv2 = 23'b00001110100110001000110;
12'b111100100001: finv2 = 23'b00001110100001110010101;
12'b111100100010: finv2 = 23'b00001110011101011100101;
12'b111100100011: finv2 = 23'b00001110011001000110101;
12'b111100100100: finv2 = 23'b00001110010100110000110;
12'b111100100101: finv2 = 23'b00001110010000011011001;
12'b111100100110: finv2 = 23'b00001110001100000101100;
12'b111100100111: finv2 = 23'b00001110000111101111111;
12'b111100101000: finv2 = 23'b00001110000011011010100;
12'b111100101001: finv2 = 23'b00001101111111000101010;
12'b111100101010: finv2 = 23'b00001101111010110000000;
12'b111100101011: finv2 = 23'b00001101110110011010111;
12'b111100101100: finv2 = 23'b00001101110010000101111;
12'b111100101101: finv2 = 23'b00001101101101110001000;
12'b111100101110: finv2 = 23'b00001101101001011100001;
12'b111100101111: finv2 = 23'b00001101100101000111100;
12'b111100110000: finv2 = 23'b00001101100000110010111;
12'b111100110001: finv2 = 23'b00001101011100011110011;
12'b111100110010: finv2 = 23'b00001101011000001010000;
12'b111100110011: finv2 = 23'b00001101010011110101110;
12'b111100110100: finv2 = 23'b00001101001111100001101;
12'b111100110101: finv2 = 23'b00001101001011001101100;
12'b111100110110: finv2 = 23'b00001101000110111001101;
12'b111100110111: finv2 = 23'b00001101000010100101110;
12'b111100111000: finv2 = 23'b00001100111110010010000;
12'b111100111001: finv2 = 23'b00001100111001111110010;
12'b111100111010: finv2 = 23'b00001100110101101010110;
12'b111100111011: finv2 = 23'b00001100110001010111010;
12'b111100111100: finv2 = 23'b00001100101101000100000;
12'b111100111101: finv2 = 23'b00001100101000110000110;
12'b111100111110: finv2 = 23'b00001100100100011101101;
12'b111100111111: finv2 = 23'b00001100100000001010100;
12'b111101000000: finv2 = 23'b00001100011011110111101;
12'b111101000001: finv2 = 23'b00001100010111100100110;
12'b111101000010: finv2 = 23'b00001100010011010010001;
12'b111101000011: finv2 = 23'b00001100001110111111100;
12'b111101000100: finv2 = 23'b00001100001010101101000;
12'b111101000101: finv2 = 23'b00001100000110011010100;
12'b111101000110: finv2 = 23'b00001100000010001000010;
12'b111101000111: finv2 = 23'b00001011111101110110000;
12'b111101001000: finv2 = 23'b00001011111001100011111;
12'b111101001001: finv2 = 23'b00001011110101010001111;
12'b111101001010: finv2 = 23'b00001011110001000000000;
12'b111101001011: finv2 = 23'b00001011101100101110010;
12'b111101001100: finv2 = 23'b00001011101000011100100;
12'b111101001101: finv2 = 23'b00001011100100001010111;
12'b111101001110: finv2 = 23'b00001011011111111001011;
12'b111101001111: finv2 = 23'b00001011011011101000000;
12'b111101010000: finv2 = 23'b00001011010111010110110;
12'b111101010001: finv2 = 23'b00001011010011000101100;
12'b111101010010: finv2 = 23'b00001011001110110100100;
12'b111101010011: finv2 = 23'b00001011001010100011100;
12'b111101010100: finv2 = 23'b00001011000110010010101;
12'b111101010101: finv2 = 23'b00001011000010000001111;
12'b111101010110: finv2 = 23'b00001010111101110001001;
12'b111101010111: finv2 = 23'b00001010111001100000101;
12'b111101011000: finv2 = 23'b00001010110101010000001;
12'b111101011001: finv2 = 23'b00001010110000111111110;
12'b111101011010: finv2 = 23'b00001010101100101111100;
12'b111101011011: finv2 = 23'b00001010101000011111011;
12'b111101011100: finv2 = 23'b00001010100100001111010;
12'b111101011101: finv2 = 23'b00001010011111111111010;
12'b111101011110: finv2 = 23'b00001010011011101111100;
12'b111101011111: finv2 = 23'b00001010010111011111110;
12'b111101100000: finv2 = 23'b00001010010011010000000;
12'b111101100001: finv2 = 23'b00001010001111000000100;
12'b111101100010: finv2 = 23'b00001010001010110001000;
12'b111101100011: finv2 = 23'b00001010000110100001101;
12'b111101100100: finv2 = 23'b00001010000010010010011;
12'b111101100101: finv2 = 23'b00001001111110000011010;
12'b111101100110: finv2 = 23'b00001001111001110100010;
12'b111101100111: finv2 = 23'b00001001110101100101010;
12'b111101101000: finv2 = 23'b00001001110001010110011;
12'b111101101001: finv2 = 23'b00001001101101000111101;
12'b111101101010: finv2 = 23'b00001001101000111001000;
12'b111101101011: finv2 = 23'b00001001100100101010100;
12'b111101101100: finv2 = 23'b00001001100000011100000;
12'b111101101101: finv2 = 23'b00001001011100001101110;
12'b111101101110: finv2 = 23'b00001001010111111111100;
12'b111101101111: finv2 = 23'b00001001010011110001011;
12'b111101110000: finv2 = 23'b00001001001111100011010;
12'b111101110001: finv2 = 23'b00001001001011010101011;
12'b111101110010: finv2 = 23'b00001001000111000111100;
12'b111101110011: finv2 = 23'b00001001000010111001110;
12'b111101110100: finv2 = 23'b00001000111110101100001;
12'b111101110101: finv2 = 23'b00001000111010011110101;
12'b111101110110: finv2 = 23'b00001000110110010001001;
12'b111101110111: finv2 = 23'b00001000110010000011111;
12'b111101111000: finv2 = 23'b00001000101101110110101;
12'b111101111001: finv2 = 23'b00001000101001101001100;
12'b111101111010: finv2 = 23'b00001000100101011100011;
12'b111101111011: finv2 = 23'b00001000100001001111100;
12'b111101111100: finv2 = 23'b00001000011101000010101;
12'b111101111101: finv2 = 23'b00001000011000110101111;
12'b111101111110: finv2 = 23'b00001000010100101001010;
12'b111101111111: finv2 = 23'b00001000010000011100110;
12'b111110000000: finv2 = 23'b00001000001100010000011;
12'b111110000001: finv2 = 23'b00001000001000000100000;
12'b111110000010: finv2 = 23'b00001000000011110111110;
12'b111110000011: finv2 = 23'b00000111111111101011101;
12'b111110000100: finv2 = 23'b00000111111011011111101;
12'b111110000101: finv2 = 23'b00000111110111010011101;
12'b111110000110: finv2 = 23'b00000111110011000111110;
12'b111110000111: finv2 = 23'b00000111101110111100001;
12'b111110001000: finv2 = 23'b00000111101010110000011;
12'b111110001001: finv2 = 23'b00000111100110100100111;
12'b111110001010: finv2 = 23'b00000111100010011001100;
12'b111110001011: finv2 = 23'b00000111011110001110001;
12'b111110001100: finv2 = 23'b00000111011010000010111;
12'b111110001101: finv2 = 23'b00000111010101110111110;
12'b111110001110: finv2 = 23'b00000111010001101100110;
12'b111110001111: finv2 = 23'b00000111001101100001110;
12'b111110010000: finv2 = 23'b00000111001001010110111;
12'b111110010001: finv2 = 23'b00000111000101001100001;
12'b111110010010: finv2 = 23'b00000111000001000001100;
12'b111110010011: finv2 = 23'b00000110111100110111000;
12'b111110010100: finv2 = 23'b00000110111000101100100;
12'b111110010101: finv2 = 23'b00000110110100100010001;
12'b111110010110: finv2 = 23'b00000110110000010111111;
12'b111110010111: finv2 = 23'b00000110101100001101110;
12'b111110011000: finv2 = 23'b00000110101000000011110;
12'b111110011001: finv2 = 23'b00000110100011111001110;
12'b111110011010: finv2 = 23'b00000110011111101111111;
12'b111110011011: finv2 = 23'b00000110011011100110001;
12'b111110011100: finv2 = 23'b00000110010111011100100;
12'b111110011101: finv2 = 23'b00000110010011010011000;
12'b111110011110: finv2 = 23'b00000110001111001001100;
12'b111110011111: finv2 = 23'b00000110001011000000001;
12'b111110100000: finv2 = 23'b00000110000110110110111;
12'b111110100001: finv2 = 23'b00000110000010101101101;
12'b111110100010: finv2 = 23'b00000101111110100100101;
12'b111110100011: finv2 = 23'b00000101111010011011101;
12'b111110100100: finv2 = 23'b00000101110110010010110;
12'b111110100101: finv2 = 23'b00000101110010001010000;
12'b111110100110: finv2 = 23'b00000101101110000001011;
12'b111110100111: finv2 = 23'b00000101101001111000110;
12'b111110101000: finv2 = 23'b00000101100101110000010;
12'b111110101001: finv2 = 23'b00000101100001100111111;
12'b111110101010: finv2 = 23'b00000101011101011111101;
12'b111110101011: finv2 = 23'b00000101011001010111011;
12'b111110101100: finv2 = 23'b00000101010101001111011;
12'b111110101101: finv2 = 23'b00000101010001000111011;
12'b111110101110: finv2 = 23'b00000101001100111111100;
12'b111110101111: finv2 = 23'b00000101001000110111101;
12'b111110110000: finv2 = 23'b00000101000100110000000;
12'b111110110001: finv2 = 23'b00000101000000101000011;
12'b111110110010: finv2 = 23'b00000100111100100000111;
12'b111110110011: finv2 = 23'b00000100111000011001100;
12'b111110110100: finv2 = 23'b00000100110100010010001;
12'b111110110101: finv2 = 23'b00000100110000001010111;
12'b111110110110: finv2 = 23'b00000100101100000011111;
12'b111110110111: finv2 = 23'b00000100100111111100110;
12'b111110111000: finv2 = 23'b00000100100011110101111;
12'b111110111001: finv2 = 23'b00000100011111101111000;
12'b111110111010: finv2 = 23'b00000100011011101000011;
12'b111110111011: finv2 = 23'b00000100010111100001110;
12'b111110111100: finv2 = 23'b00000100010011011011001;
12'b111110111101: finv2 = 23'b00000100001111010100110;
12'b111110111110: finv2 = 23'b00000100001011001110011;
12'b111110111111: finv2 = 23'b00000100000111001000001;
12'b111111000000: finv2 = 23'b00000100000011000010000;
12'b111111000001: finv2 = 23'b00000011111110111100000;
12'b111111000010: finv2 = 23'b00000011111010110110000;
12'b111111000011: finv2 = 23'b00000011110110110000001;
12'b111111000100: finv2 = 23'b00000011110010101010011;
12'b111111000101: finv2 = 23'b00000011101110100100110;
12'b111111000110: finv2 = 23'b00000011101010011111010;
12'b111111000111: finv2 = 23'b00000011100110011001110;
12'b111111001000: finv2 = 23'b00000011100010010100011;
12'b111111001001: finv2 = 23'b00000011011110001111001;
12'b111111001010: finv2 = 23'b00000011011010001001111;
12'b111111001011: finv2 = 23'b00000011010110000100111;
12'b111111001100: finv2 = 23'b00000011010001111111111;
12'b111111001101: finv2 = 23'b00000011001101111011000;
12'b111111001110: finv2 = 23'b00000011001001110110001;
12'b111111001111: finv2 = 23'b00000011000101110001100;
12'b111111010000: finv2 = 23'b00000011000001101100111;
12'b111111010001: finv2 = 23'b00000010111101101000011;
12'b111111010010: finv2 = 23'b00000010111001100011111;
12'b111111010011: finv2 = 23'b00000010110101011111101;
12'b111111010100: finv2 = 23'b00000010110001011011011;
12'b111111010101: finv2 = 23'b00000010101101010111010;
12'b111111010110: finv2 = 23'b00000010101001010011010;
12'b111111010111: finv2 = 23'b00000010100101001111011;
12'b111111011000: finv2 = 23'b00000010100001001011100;
12'b111111011001: finv2 = 23'b00000010011101000111110;
12'b111111011010: finv2 = 23'b00000010011001000100001;
12'b111111011011: finv2 = 23'b00000010010101000000100;
12'b111111011100: finv2 = 23'b00000010010000111101001;
12'b111111011101: finv2 = 23'b00000010001100111001110;
12'b111111011110: finv2 = 23'b00000010001000110110100;
12'b111111011111: finv2 = 23'b00000010000100110011011;
12'b111111100000: finv2 = 23'b00000010000000110000010;
12'b111111100001: finv2 = 23'b00000001111100101101010;
12'b111111100010: finv2 = 23'b00000001111000101010011;
12'b111111100011: finv2 = 23'b00000001110100100111101;
12'b111111100100: finv2 = 23'b00000001110000100100111;
12'b111111100101: finv2 = 23'b00000001101100100010011;
12'b111111100110: finv2 = 23'b00000001101000011111111;
12'b111111100111: finv2 = 23'b00000001100100011101011;
12'b111111101000: finv2 = 23'b00000001100000011011001;
12'b111111101001: finv2 = 23'b00000001011100011000111;
12'b111111101010: finv2 = 23'b00000001011000010110110;
12'b111111101011: finv2 = 23'b00000001010100010100110;
12'b111111101100: finv2 = 23'b00000001010000010010110;
12'b111111101101: finv2 = 23'b00000001001100010001000;
12'b111111101110: finv2 = 23'b00000001001000001111010;
12'b111111101111: finv2 = 23'b00000001000100001101101;
12'b111111110000: finv2 = 23'b00000001000000001100000;
12'b111111110001: finv2 = 23'b00000000111100001010101;
12'b111111110010: finv2 = 23'b00000000111000001001010;
12'b111111110011: finv2 = 23'b00000000110100001000000;
12'b111111110100: finv2 = 23'b00000000110000000110110;
12'b111111110101: finv2 = 23'b00000000101100000101101;
12'b111111110110: finv2 = 23'b00000000101000000100110;
12'b111111110111: finv2 = 23'b00000000100100000011110;
12'b111111111000: finv2 = 23'b00000000100000000011000;
12'b111111111001: finv2 = 23'b00000000011100000010010;
12'b111111111010: finv2 = 23'b00000000011000000001110;
12'b111111111011: finv2 = 23'b00000000010100000001001;
12'b111111111100: finv2 = 23'b00000000010000000000110;
12'b111111111101: finv2 = 23'b00000000001100000000011;
12'b111111111110: finv2 = 23'b00000000001000000000010;
12'b111111111111: finv2 = 23'b00000000000100000000000;

     endcase
    end
  endfunction

  wire [22:0] m2;
  assign m2 = x2[22:0];

  assign y1 = {1'b1, finv1(m2[22:11])};
  assign y2 = {1'b1, finv2(m2[22:11])};

endmodule

`default_nettype wire
