`default_nettype none

module itof(
  input wire [31:0] i,
  output wire [31:0] f );

  wire s;
  wire [7:0] e;
  wire [22:0] m;

  assign s = i[31:31];

  wire [32:0] p33;
  wire [31:0] p32, p;
  assign p33 = {1'b0, ~i} + 33'b1;
  assign p32 = (s) ? p33[31:0] : i;

  assign p = (p32[30:30]) ? p32 + {25'b0, p32[6:6], 6'b0} :
             (p32[29:29]) ? p32 + {26'b0, p32[5:5], 5'b0} :
             (p32[28:28]) ? p32 + {27'b0, p32[4:4], 4'b0} :
             (p32[27:27]) ? p32 + {28'b0, p32[3:3], 3'b0} :
             (p32[26:26]) ? p32 + {29'b0, p32[2:2], 2'b0} :
             (p32[25:25]) ? p32 + {30'b0, p32[1:1], 1'b0} :
             (p32[24:24]) ? p32 + {31'b0, p32[0:0]} : p32;

  assign e = (p[31:31]) ? 8'b10011110 :
             (p[30:30]) ? 8'b10011101 :
             (p[29:29]) ? 8'b10011100 :
             (p[28:28]) ? 8'b10011011 :
             (p[27:27]) ? 8'b10011010 :
             (p[26:26]) ? 8'b10011001 :
             (p[25:25]) ? 8'b10011000 :
             (p[24:24]) ? 8'b10010111 :
             (p[23:23]) ? 8'b10010110 :
             (p[22:22]) ? 8'b10010101 :
             (p[21:21]) ? 8'b10010100 :
             (p[20:20]) ? 8'b10010011 :
             (p[19:19]) ? 8'b10010010 :
             (p[18:18]) ? 8'b10010001 :
             (p[17:17]) ? 8'b10010000 :
             (p[16:16]) ? 8'b10001111 :
             (p[15:15]) ? 8'b10001110 :
             (p[14:14]) ? 8'b10001101 :
             (p[13:13]) ? 8'b10001100 :
             (p[12:12]) ? 8'b10001011 :
             (p[11:11]) ? 8'b10001010 :
             (p[10:10]) ? 8'b10001001 :
             (p[ 9: 9]) ? 8'b10001000 :
             (p[ 8: 8]) ? 8'b10000111 :
             (p[ 7: 7]) ? 8'b10000110 :
             (p[ 6: 6]) ? 8'b10000101 :
             (p[ 5: 5]) ? 8'b10000100 :
             (p[ 4: 4]) ? 8'b10000011 :
             (p[ 3: 3]) ? 8'b10000010 :
             (p[ 2: 2]) ? 8'b10000001 :
             (p[ 1: 1]) ? 8'b10000000 :
             (p[ 0: 0]) ? 8'b01111111 : 8'b00000000;

  assign m = (p[31:31]) ? p[30:8] :
             (p[30:30]) ? p[29:7] :
             (p[29:29]) ? p[28:6] :
             (p[28:28]) ? p[27:5] :
             (p[27:27]) ? p[26:4] :
             (p[26:26]) ? p[25:3] :
             (p[25:25]) ? p[24:2] :
             (p[24:24]) ? p[23:1] :
             (p[23:23]) ? p[22:0] :
             (p[22:22]) ? {p[21:0], 1'b0} :
             (p[21:21]) ? {p[20:0], 2'b0} :
             (p[20:20]) ? {p[19:0], 3'b0} :
             (p[19:19]) ? {p[18:0], 4'b0} :
             (p[18:18]) ? {p[17:0], 5'b0} :
             (p[17:17]) ? {p[16:0], 6'b0} :
             (p[16:16]) ? {p[15:0], 7'b0} :
             (p[15:15]) ? {p[14:0], 8'b0} :
             (p[14:14]) ? {p[13:0], 9'b0} :
             (p[13:13]) ? {p[12:0], 10'b0} :
             (p[12:12]) ? {p[11:0], 11'b0} :
             (p[11:11]) ? {p[10:0], 12'b0} :
             (p[10:10]) ? {p[9:0], 13'b0} :
             (p[ 9: 9]) ? {p[8:0], 14'b0} :
             (p[ 8: 8]) ? {p[7:0], 15'b0} :
             (p[ 7: 7]) ? {p[6:0], 16'b0} :
             (p[ 6: 6]) ? {p[5:0], 17'b0} :
             (p[ 5: 5]) ? {p[4:0], 18'b0} :
             (p[ 4: 4]) ? {p[3:0], 19'b0} :
             (p[ 3: 3]) ? {p[2:0], 20'b0} :
             (p[ 2: 2]) ? {p[1:0], 21'b0} :
             (p[ 1: 1]) ? {p[0:0], 22'b0} :
             (p[ 0: 0]) ? 23'b0 : 23'b0;

assign f = {s, e, m};

endmodule

`default_nettype wire
